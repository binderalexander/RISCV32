
module riscv_simulation (
	leds_export);	

	output	[7:0]	leds_export;
endmodule
