// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:40:51 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SGam8xW6TRBYQzdjXPTgG+iu91+BVR8GmH7/m1fPm+p7MxF23lNdkPCrqIpb4Wil
ewVpITZ4RgE7f62WK2PdxA56svnV0588djhOaq9zIryFEnPml/F5h66dQXUe50Ky
dCYOon8Gjy6FA1tyasrNyGiZRlI/35/ehyu8/NBwwrU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 68208)
oW3+cqjX3+c6nKSWQuP7pGojtn2dCv5rUS7xWhuIcVJU3w53hXvdNLJCUW7TP/QB
oZgPlpu1kTYdsFy56x3n0tdYmPs4vcHdmP4GKvl2SkolOIlFLpAvw5J30bPwP3mf
Byi21b6jBomJHyDuCmUgRBUJmA2hZC7VYsEEqm8D7JrupKr6wZ0VpCNWxKCpJDtX
riWJwg4jOLtm8RaO8tapG2blsN/jQ3x17NTjfIXDmLPpiN/HTVuQTbJdIrxO0q2M
bbNjaGuosXaC2UP/2hbpcazRXymTcAzSbf94yxHPMqYgABVCU2FYGvRwiTwzCf+b
Y6hnpLD/6hK3A9BTdVJaSX+RP1XuJ9OaQtpzKfXs4Djtmqw0Dhkxp/ARqKYg4610
P1iJnsSOeGiBl3Yh75SVOd8WtVljChw4XqTZL+09P7jZqqhA+A4tAvFPBMONKknd
oE1WPqExNJb0y8NTRY+m0Zg3Rw0qnfeBH+r8983ALbkS9+zsV1xcqaGYvp5MRl1D
plXXHQUwkkgZzO00YsHfVXiii2djZvNuo12y3eJ2BbO5trvAWKdv/qjetO97WOkB
aQOpuedx3hbHejSMN1batQHR7ku0WlJokXV4IyjrRdsYM6FMbqQbt5ltXbVxa8T0
2Hv/Z6kYbJcVntIvYCAfbDBUgWdK1+5CKB61uF6Ai3bj3qN0vnuUezCni4bq88yM
ODsd+pLOnH/YTDDqPYghpkFx1lCRKQGXK3rBBGkAOh3rSE+RPIaYMB/yF/6TqP5j
1dKtLeUp6xknemGJhNv1w1wKt2S3OKc9SrwqBWDUqRUnBXadlTSCaEzaJZrkN3d9
J2LBEmGFMQhBoa9SbR7k5yVS2pS5ZBUc/nbGiJCqSmBxleES0XcGXerqRL9AUtHS
9jaED8jF5l1DRbWnHku59NX3SWhPV4SkAVxWLZmUF3bI+NPixvu/L6tWbF0fi1kO
mJFT6XrBhLHfGyf63YsNbWZzgqOUjitrbH70etJ36yO6Xolhj8XOPoOrYtyketQ9
G8QOhexNovCJjUHAcaPFKHpvrJ1RSsbR3R6jMRG9CBZW7t3DiyPgEPR3Nypr4+IV
jGv4iWmM/EoA+VZO/+DyLL9AXwybUiH4G3TjQjJSWfmFkzh7z1vPczJOGWNlBI+a
9S6O/bv+h3bxFto1q/Vxd6eIGMGMAAk1CIHXdaXS8M4bwOi/Gr0IqJmOobrBtU3Z
foTTmOPUGPiokbtuHlgCClMCBHUd3y1Sp6ZJFW1JzJsCJgumq3XPUdFt97NEoJGC
qB8R4F2pjLoPT9PEecuJQe2rpqvShMo4EFqyLAMutYJLW0yRl0JhJ/CuZRuQDC2u
A1wjrStVMNtEF1rS2gLLX4s+oyS1cXgTZS8PHsK/saLj+xIQQUTi1nGVFBgRnjD7
YeXTPfO77wSAuPJh46kY/htTSkWMbi0QHNX+1RGdyJK/jEOjmD2G8WOgw0A94bmo
3SnHvvIr1nStnoqlhY7iMgkWZbj3mtoKGCJL2756lY7POaV48zvOzGb2D0RSmzN/
1b1QFiscPrv/vuwmGVehZyCffuvpNxLjwx114LLZupE1q3yGb9DQ+qrpSWr/5nTS
RoYKgSsAWAqvrQlv6zYMFm5QQbmZFETb3RLZREsyHcffwkaMjXHRwsEDTKvAs1hf
gG+C3mcchgfxQp8sj6rawWVMl9jmhJjii1ngHMcPaNaeaSxRIVLpP+C56lR4eQu6
4dzRtOsarGVO8L6udhh8DkU5sLUzFb/9SrKIxgyv05nov87/XF80Bz7o6lgvRNkT
sYh1xu1PvG64E/kDnb9XmWhSfIPJPPZ2w5FnNxgfmU+FgPRlclvEtHhnTN38KERS
TY+wXn3EZN2Pz8baLW7K1fFUtKRVTGE5gvNp76AQ5hWvYz+AvngE+omr89chZ+fT
lwkfKb+TOlCHBtyDJjVTU13dw9bBwQZSW9CrcoQzKLCvU14GzCgH+zQIsWOzT9YY
Uw++4+R9S5hGr4n5Uij76Kpna8dp8jRM3i5IwwxUdJeAxIPCiwb0L4CgZU0u65EA
fjuVTYm0nOXDRre04+fIhRkq/d882szhAS/fNr+TX692h5zn3GFd5pCmjEBb73hr
YxlngvsYLmtj0RMuWAUo79SlsfwJ3lBebfjLlhvs3mH/9sY79BKslArR6C8nCXUw
AhY4O3KpTmZyfkASHxojUP2WaU0AXwC1CyYRDccDWCJNil7M+czNwOMGEhQNsoDh
WNjE7YU8R9fiMQPkMyCXyg2Slwk9kBLza1kA05yHpElq8UnB6PhOWhtxYI/DWOMX
97UAO58UKLYJcsawnOhRKAnympnDhl7szKxTdCOr6uwPvbwVxJu6zxRS2U5/UAkC
3tSlwwhJEqGaAN9ftDxW5fswNWV3jtrXwldVIsVUM3EVVc3ETeFL4z5GTIxEqZgv
QzpCI1ZXrwytK9wqBKJpv8A0JJWwmTCr74a26ELpNWn+GMxAxVDsoOLgbxuhY1Fs
yQo0aAV0broDl9oEdk0Iuxspiuqu8iSarWEwlX4ILrMBxrpu0jrVHLMmHEu/gtOO
tU1G4UNKwORju+rVsTx6a/H/p68UgCyXq6HZ9k0c8zbCPGlrXk5Vd/+gCKSgQ+LG
ZhOz8BjfhJq4JdCi7ZIfcCVM8+CIHSLp1QJ38JSfKq4rlpKEEWyaF+9to8+Xf1N/
r4flePV6/9QnlcHEgHRwSONhR0RijtkV4yOmhwvVkcRjaonvOfWH+fpd6eNpglz0
ZjUXKnqfKEmZ2+ayqpD2iyj9Dsp1qfpkaEYj24UDAHUusI5bgQiw/+Z1hr3FXLqn
peNm9zzerL7IEErEJUDMERNZJIp7W83OHVLysOUrJ+yb7jCmL8DOanYG7Gco8Slw
WvP6ot1K3KNNWpUXupvnRmmcFS6bzjgaKB8uzrPO1D0UKqaI/t0MTbb+rJMR3v9B
YhZ3m6BqiMHvhePv1UJjWYAgtxHsHCDuoWVzbQ5nyMNZTMpp639UzrSip4QgfLQE
VA1ChsAYp1H0Je9UGoFOn7WbqDALotWIzf0U11X0mAsIpuum5lTghU7b8GBBFydd
hnmawl4p+FQ8N6odH8bDvvj7XkpDb7iGlzVcPYhcEHDsM+fyLnWml2ALt8PzczNF
mocMY60kafaurFEaMVDtXlotBQeMdj1uvr1Fhwj6YoN0jDQVT7YRJRINjy6wCu+J
4q4AkBZunvzaUPChHvBebF1h8dECbF+Gd8oRZW97Qi6yl//taCJBhYFXT8ho12S6
O9N/8pk95BAOHZ2HFyUFfJTyqOjhuBVRrcRTaBEJ9Z6iY6+t+bzcR374xmmmvQT2
05kPfYaiEcovy4wOYq0YZt56XsIAfpLQgYVSE0bIEB3tNAja7RWAYyyhQy8FKzB7
t2Uvphlv+lqS3eYp+QC2e0SA8NI1eJ0qlrm5ZkGjKyS+sPh7KD2oKa/kTWmR2z4S
A668fOh5OgPek1dat4vsznRGDCaDqK1+A546BWdzC4QbEMtHInVjf0WgSqn76lpZ
5rIxXK+Oy/4DfsfePBCP7qaFFr0zZ6EkvkoYV4ZDIyMzykwRp2PNQ+tGFZu11+jX
SJLADRxet2DddYeepFYzH20TvI4F9fYgLptIYtTUtt8SWCHYTgYRCqAuTepMpEpf
jEEDPQJjukepyjuKMPN79JON6RS2w5ACng6gZUxT1013PWSNliuPI9GTL8Qr90Yu
VphxxQ1dmqOD0ewbwaHVuUVACtFQvLLoGovzd6fubfVI5xvf7savGYZehak8PPyR
d7OBVtfg7/59fT3PAQED4uMKKkgXS7oAYB8DHq4KGpafkvZs+XoeDfuTNekYBOHy
LAAkUu0HplZeHNV/tP+8CXZFAB8hszmPx6Lf7IN3FQqVnriBQcZQJ4tY6CHG/yn4
u2XisFTGKIfcDs4zcNTYKfIBDi1vBqy3Pa/7uBZ9rz0utTYHcuvXkR+T9+hmEWBC
7W6tE/00woH911eYLdraETgCAUv7lJ5IlM8TBr2GbmnuzSEsEceleGBEvaydZYvH
ygKxmzXxsb4ZnFv7pzIx0PaQo6vPzeXSTmCY67jy80cLheDIUFjKpzvsdFCLrFk/
GkWnXOAWh34mKSLmQNhGFxgXaqAMApgG0SONY9ksdD8vDEJee8CIcUoA080CYeBX
NRuBbTSajyhSCS4BMCegJg0sVJU7WYJF+FTPk+WnzYXM4MRkVwXqBRLBywODBPm+
5eXBMUyMo1+mELFf3a2vyJw5Nn4IsPkGrHGLU6inTzclv4QV+vVmqI80MwHuHGob
Bm75NDtucHNpfnSUkt/3wkGBAFkajabRPqhKnyKjHx7WoEFZeU66OI+866fXsLwP
cbMX/yWv4Cq1xdtHAmtPFVfMyD2GPkUvXzeegSF9lyElSqWyVVk4wwfRdBJfZ3yh
U94Xtr2O7kxMs2Dr0twhawbktbRsz4egzLYmoorC5pOqDPUnp7Sv+T964DrVZv5T
RC6aLrRVftzAe88MLpm802I2+KIvu4w22yR8I8xPraAV5zkMZiIRxkHiw/Hm29pp
+F9YtzAPfwwi/QlrUUyCnfiCtlxZK7W8xYCxK/VSkqozZXsfzrCBpV+7st2Bo6q4
GWv82vkfE2+UWZw2KiA/FlQbo0QQl0NwdGtHu/h5//bxVpp/3FClFqiztqu2iPdV
sO+Ab18thxRQJlnvH5odPGKGQqQdr2I098t0SvdHXN7X3xpM+8/ma4jvwP6gGYEk
QKEYJ92Y1T8GDOPlkbtEEc249uhtqyDuuWHzixpYjAiLbOM0vvOLLwBEWFFsqqPI
2T5e1wBpYRm7Bt4rn9QSvZqf9+ZPjRimONYZtR82s00bQ33v6vmZH2+8IoFme4Ce
m8wgRSaHpx8pCZ8dHOjZSuTC5SY2sJaErIj1nKzVM/c17nZjsveUREYbtMTyDat+
wsrdJD6OvryFx/QWilB0JY7Vlview9N3uWy63po9dFqdNkNUcmP4NeaPAI5TuosM
FiPv26p4G/D3SX3NU4xOElXcuqiFER8JT6jgGqGFSaM+ZbQ32IN4QKJKhBwwau0e
OGy2RQ35TSByrkgGSn5+37ZPtztHLP6xMd2n3axeN11hN0aLRh65KRYrVDuIDKxi
/7ovk8pywBMM/Y7G3imRdGUOrcRvjKJG58KX5hcs9VapdXE3udTB1BaTQaLEsPZ3
EmZFGs3xW07dNtCtGkE/FGdGNMJ01Wfv1uG5rDmfAQjjM95a/2Z6QyAIwlCxL7er
Kmmtkx5BxavRIeU2OpUYj39CGCsqaxJNl0mxSpUL6K6Ee3OgaOKd8UKj6gW2PNNK
xGTdIHdcOXYe41ZDtasISezS138rF+oweuy6MlMLiOKAqInSvpDx/WcP8Ii6Hkko
J6UOkDbqkylzU0nZZ/4ObyHhzftyQGh2ndiy9viceH6PD+PpIf3k0+N5SP3w4DUe
Ag/laLgCv0wMc5Y2gJ0H2GDPUVvlUFQcIWvM0dYbcFdZJ/sMVnnnXtYwv93YLEoV
mO0irByYzufx3qviKeex7KFcFSXpHRbYboekPg+KqRyKV/vECGrgy/EOorGBbCTr
l4xOLXIMRxfKMWUnniGxhOqDW9Z0mYGk2vBgwgWdvk8yjoNiH2Ttssdg5aVyCT8Y
k1bymYwuRXG5OaBK+U4d0R8BYKrkQWm/RDOD4wnXuhofUeJpfUQgapt9LNorNruY
snqNhNH3mEbewnWQ8Chvd5me2+kjX7s/XKOJwgvpjByCWG8YnsJNMQOaRygaKOyN
Oz0Wa9/6TK0mM7kq0IvLJ6QngDlZxNeloEUu38nVUfMuS+i0ZqFRBu4zG46Jep1z
LuQy04coV4XxY8Qv0dCjVLM8OtdlixTcQypCeYqG1DWE/zcBuSwcArS6KOxNn2/y
eZdAv+S3hbrTeIympwRfbqahkS0kOLxIk3bRmLjtEjZg1pnwVmYcqSwlNbz/8brn
rNCHRNtGz1OuailPuXcfjMLxs4gujDpltoo4e7RVb18RydYYLbyMV5hr0a/XgW+i
QenCUvEWnKQDyVD0ENkvjus6i5QpStO6gXXgWgVYMhr3vooycHUcdC49obOQMwHq
MFL8QN2ofC5cWAKCHuICUBCuIIl1U4yu8S8fKJ27D5bYmMrfGxhF1f/lzKeQJuBL
KJRzyvdyCx3Sed2qBc9B113pjkvjI5VxbxlDMvyk/5oZmTOS3ysLRMMT41vtN6jB
+9HhIYx8pQPXc59oZF6a/J2sdBSWvBVzdolJAqGqx+9xCx5nspGG0DHn0R/o78Ia
e8GPUXZf7FnLmi+0kUbLr+V4ItvJ+2i7uCilVnkraB00UZ/rE9VnBuAeu13JdpNL
sOUvGvifMFHrgIsvqi1wBAef//L72XcNWfzgG34V3l4GHs43UEhIQslCdlgaHtLc
K9imaZbaTR983dKS922Ln9dUVZSCWhL8V19CqRxVEnW893m0WB2fo9mIo/Vr2QgH
aeR5ME+TRzeFPKKT5a7mXBerWqLOWXWkUbYlt8sgpYH8AzC0Jom6JMdzUmXDmPsW
3m9zgGOsEgijH8022c3sBimBX0+lu/xEdEkj2KOKazeXscanKTvmleBvWjBk4+k7
RCo5HjWQPebInENlCZ4kRe3S8W0NCH75iSWHLMLCzQe04jBEu2MjZlVSxl0u3XSI
8HRMi2OqDLP6tYqDz84hFkxtG6hJMvWuej7JiNrfC2KeLXAnp/w0bsQlxURGLWgA
gP9eC7wyztg9mLCzPXWfT9OcwHgsjiUBMlClxkf+lrT9wbOOkmRJlbc5BAdBW01b
BBtS7NPuZ8WRy6JqQpoA1P0s67iHHWKCqxEUCR8gZoey01fsXENHJuwp+5cviMaf
JxF0GWmw+xKV0yzzo28QMhEL2h4A65Jbiw7gfj+g0vsTqLf+kzE8MfP8y+OhUlnZ
v6lnx1F+1lfm9LqOiBdekRJKSNXIi2OLpBMGCcFUA7EVNNRBQsXSUA6tPKqka+9X
0741vekvU2hFNnuS53csphuPPUyd4PX/fhefR0jTlYd9OXdY/fVH3DxETqcYYXkd
mf9tzNS3xKNRUnIBj4o2cYV3GS5bsymgUg5fwQffLFv5sgJ5bFCtXwYvqi+L2T+p
RTq8UB/Qz7zPy2n28LrZ8g1LlgalF+SyfobGvwuxEDnJ6jfNlg8i+gopXV6u9kac
xcNeztCqjQW30qGKGXWqOrUd1Jmk8vHpm22GVq4vxT9ELn7Eydbhjqa13BMFjniy
O/yQ7tZVyijjI3NE08TO3x67FppSGGrG9lDnZrQg24rLi3z5KYlmK/lEdDlJRWFy
1rbGj4YQolfkiTANIhKanuBrLY3aN+7EKbU0wTxQldX2ljaqS4CtUEKupDjKgYCu
VxYDcgBKg+uMQjpIOs8C8NIrlrDF6Mu2SxEjllKKU4A2zXDR6FJpspetHto+RLxg
N1DykjEUXdMwgXekLEoN507QAbx1WJVmoXwocCajCMFysUBmFYcqHmc9ZfuKLxY8
0Em/BlJvoO+KUe3OXRMx5bghHAFLJGbR7tEuGCVIygnH4WI18rFZk2OeAAq/9GdL
gXS7t3k8Ki+aKv+bv8uueIvMr4yKIKOTCk7fACE/El/q8ebi5BT4qFB4DKg4cmhr
UeJAeJlSRfUpBYiU/zK2UymKg2Vok+VnSWMmBYJdYc/eMZAxmnQNDYxYq6vAMj/X
STgQugzTAV3HqCj2v30AuGEoWhETMT9JBzZXWH4bj7dunQrmjk6o90I8DpwSyQZ5
rCE3OoutjcgdUIZ1E4oedoArsL2pCfaclPYsH+n8x1X+QWxCi7xgUsX9DMzfY8pM
Qv9rhiV1GqcO6mGzXCl5YgZktAdzpnRs7WFtDTcWUUSh123e/257z+hKZtwfxCwn
4u2f3Fzdtm3ea+Tk4wE43He3nToV0bvUxUPvmFRxYoIAVxEWZ8jxcrCyxZAiTK/Z
Pr0rkBKCIjw7NWj95cJX7pvms8JM67X5NMv3aPmQaW/RfrpHHcI6KL3SQqvh7uCM
nYlGP/0yIR17sOY9oOX5uChXsqP1Dac9CaCpGkfPebCJQCE+aoQwZy1wmfXVTyMp
BubD59R1EGfvLik8fFK5eVmm4eZpUg780VLL7BYiEDEuFb2sDWuy4CtduW18Bhip
LMBoaGyxNwtRNQRLqJFxBtBWnv4Ah8XoW3UKFHDKhQ80A2TABDbmEWx3C0DEGiBJ
e2Q0iC02FxC+NWnS+1Yb6/h/TiQuksdwRaArJpeCzjMA8pfWZ15BfkPlTerGgjRx
qLJe5fyhwmwCS6ILpCcxsGsHhBHrtYBYuMMaX11loF6vCToucktjh6QgT110I0aF
o0DldiSzf05bnBqltnrHI7/UaZfOoBS02jhtQCCPL7SnWbyqyMJSYTdQ97ayrKTZ
emtwZFWI8BLqqpFToziTYuuuZhTokHaWn+68GdIp2iZ236e5ipHxZtTMxAKEPnh9
VU7dIMJ2I9T20xA6KmdBeqypRgrkJkcahg1csV2MQhZS3A3Ry0PoiVNuTmqG2zDX
tv3bGXYU5KVXbmKeGz5kaRsy7s3pwn8A9FVJhr9RQdkIuMLFsgzrbZe0yAqldWEJ
YDX5syCMv+oHuiAm5kerJm9ezbX3uFHq5PZi0cgg0bQlpF+8VsbgQkT0H8I23LJm
nMTxx6X1XohM0F+45M1Nib9kgBZENpenFY30Viw9mRVuMB0AKwROr9KIy2Z3BJeG
l5eJegA9RsvXvlbTQwDXSOLaq+q75j42bF4/7BzbePIhhkNBH5dtD1uFV5WtjKCr
6Hp/4apgUKy7ltl+XwV4VuntZtqNLxtY/tRi/oXa337H+Q1AePJlZ/5dR9SkfyoZ
dcrOrVuOH6tCIjS1JeHgW3+uadSsfxW3QGHoG8QoOoAdwmLcTytIbBSpo6o8E5o+
46mxjRjhswpU7dd94I8U4fagcPAAl1lGxnxkn1hWA3mXALIB8AfxKY5NsNA68iYQ
dSWqWjDNwr3cRJBK7Hy+wqDB+Vx3gdq8Bjej23dNPbqSVbGkPunmgo+m9ebRSfVA
aK8sU3r86OCED6/JL24mIKmiwAoOwonrGBjHHJAFCyp5v62OnEDMxqvnYnuUfT8I
Ne+BL5R36h9TxjkVYooO6I/KG5nMClSe3mM8nxgft8wSHzMaDQvUJjIjEN/cVreG
g0vzTuGUcL9Sf8DgUoUhoFPq+AmJ3kTufU/5/buR2AxH5NUoB1PxZ/7xQHsFCFgs
XjF1bO1kq2nGMgT6dFBJ/G1QCSfyVXmjDx5hOWA8vvZFlL1cCPkhUe/JJDJ7c94b
YJHMs5Hy0NwzoOn3KKh05ahSNYTMFC9tIRS9FuEizO5MgEQh6oymsyh5lOemyVAr
cXRE8R3ww/rGxAHKOePvTLvM66pKH1hOXP6lIPMV2gic8A5EatLOGcFD64KfhN7c
JdW/YW/gsFevN3jHbr9Ckq2KH9K3s4wKBEzheUrAXHy84ijxi26+WngbRpBJuoeE
0aNWkGd45OrlywwXSUTeepFGHFXVgACwBzi08+why5cbkpEzBs0exfoWqg/l5Oxu
qFDw0DQAPIGOm0cuTZdpuQdmAMwIG4oWvgmad5r1O6WDrXba482ODTfjTa+rNzGg
GJgoci6FcGmbDu/2zMq6kqer8Z5KnmUJeonWmpulfAdFOx4w1/1ttZGYBf9E5jy7
8a4hqZJQr8UmLW27vTzoQck0n8dW2uGvX5+k4stbcz6CZA0P08mmt0KwLcYPpkNh
e7aaq3n02yYkdAVpJ3rCG9MQX4atuBopfq1GQmw8eLeDMAFzxv6j9Ev3qsqinMAv
gTes8uMwPEyCAWbcQoET0qOM6ydmZbNWyMEdS43vhIq4MtooMk4wiD7RNrMz+LSn
GF9WM3O3aETa34UxNTL6kzJBeEfm7Eii1cKFlHdFv2DC4wbx1YC7+znZpYJXeahF
PdjMKAKuMJYowrYq2B9lvs1vpJs3Ofln9ERqR3y1pQGm2LIsii8Spcvwjj9+SxLT
yaP9wX5R2bDESLc3pxj4B5LwGJIlZK1P3bWVkdDD5hMGwi/DZIlDNfQYapJeISk/
FFYnSxbGkBA/Q0KVDbHiqt90n5IR5laISlaLbIb6aicjVtPCUnjX9Pf7lkxeHCkP
Mtgq/wMUcySYtcGyyHvjOHTbPxt2XjVqETH2l5Xq1weZ8sd9wyk8wAIARCAwckWI
Nhuw9NsGPQ4vvgYFjfFT5c22pH3wjYmuW8dZ4QTI9wVp3kNk2Vv5BDs/ltnK2bue
CaF3qrxYnWyx/t5CpBBxNLFTkk7oI+03FJM4adlCXnzqmgx9tbFXtR4ddXSi/7FV
fWY7YK9nTNzbE+Af7ORFUoatR0vcZ4b08NPbHEkygFzYwwJhNdnx+3UtJQe0A/Mn
597o8lijAnbB9R6QOcWG1lVMNQvqFMNBKj7cg0RNWDfTsL3ueefMIpCDMNgQiqNs
5yDzR09M6wH+2nEccaqit0jIYdg4IABeWantXJv7RYljOyId1P9yUGe+eIYOTK5v
p9AYIHq/c2S36iDp12z8Hk3JPTCddwID0Yi9q8IxBo7AFyE9vbaCTcTUIbtj9sNf
3O3VV5niwLr3fTlXziIlubZIpHITVlEqBrcIxBTvoDKQ6QYbSvuxpBTObDBbfzdw
m9CMREEao9DIyRDucDn7b64lUmzhaAiIcxA1ryb0jVZ0c0bn4BJe9+5q/9Q5wMME
uOoUBORcjOQzj++wd1mHvXd20Y9apRbMrthTVewRjcmcgr+TkCTGrOU5eWi7kY7w
FVXIh/kedSYhDH0O5EtHPRMmkCPl0vxgBlqV4MKeS1Ttrewl9ue/wPxpcPaexseO
DpsC5U3U+l75FOKEZua/jnE4AZGIVF0dJ28JbZ6epPaYhJC0A6OGplHrAzt8t49a
t9qZLapq4Ta2W5bSyBvg3HgjhhX23LRdaTkPgx7rgLdq6jA0yzibB2tutNDQUl25
nbku8LZkydqOfDZ5eM/uKSDcqQdkIgPGMxGC4OTpdjkGGmzuFAi4g9qLG6+vx1Z1
CBBqgcxVMpe+DYEkuJ4msQkue45thp1ErxLbnfRT4a0/m/OxDjz0sV1PbrgKr7gq
aBinYxRdN9Ao+BjW2jcUpdEMtNzOozlgV60wDa6yAeTCc670lzroOry3+mca3O9+
ry2fyXChYWIzWXN9vUfHJ6FiMdBBcbpnfnLv0v6UXY1GXEytEsF0LrUayyUZ/s9p
s0zVclNQaVxNPsK1YgW2JL1JpWUFi1qxaLRXqfBiuqdaDJNjm4Su7Lef4Ui765uW
1E12e3/F9FyCl25hrb8KzgoVWTO2lEyAFdu6tnbBXMaXtDCz30eRRYE1+fDeYFN2
dJzPVTU7dXw8t0/GJBloIxhGN61pOb+WQJtyDd76x1ti2QfOL8SwugdfuNFVludk
niNrjuGDmmOXrxdq61LVWf8gomOvwNeq1rMEWxm3sEJgO421yk4iET8ASFMj2eNp
OCvIrRT3P4Qst2JGbn5lNDKmwyYeYCY9EuRwY7v5b87Rd3ACO+Wg0x35+iFtukhl
tOK67gxSvNMZCPw/HIMlHWoW9HJMssSZJh/3kN4GWObDLTCPLhnppZ9dKmqYMo6t
Bbe41A+HjblQTuLr2ctqr+sRdLrM+/16A5Sr4Owy+ClfRSHM2SGWZJCQ8/59Rj6R
b95aQZxP1fTcCcos/pSFFae+bHfVWrTg3UqT2Q5uDBt0Avo+c/DYMMw2DV5RKx65
BCFDpa+RedyzY8kv4Zmi8sMOKovC/Hf6cI5N1yv6+dPbyfG33gJFKftAZ7MRidoI
L7hwy27Nc26Xd6haa3r4iQiPyFmyMVjwsOGNA7lfvZ2A07pVHzIq2EtCQlwV4HaP
IBzbCFWoB66HKVrpvbYJAoeJooBNku690iMZbTVL+/DoqmCslZdIXfn5+cBUdW/8
7C5zqsjMAZ6n0p5z4fB6d5L1s4IBjMenMpTxz3AXQkM5En3620fkpBp4CW+6MZbh
yBg1nsad88tJtX02fE7YtinW+5MuTbb+5M+0DfUGgszwRqPeDWeJWvSey2wonml3
oari3xojEOFeIsd5C0aaCVP9QhtDhhQAyL4uMy8g8zRfwC3VeSeBGCB9NYbSg66i
v5cL47D9j3nOCQ5uT2m699CLb1vo/QvQBdw7XrcJXOHQghNKdIZTNsicVqJLOyqQ
q2/4cckCy3LCMn+pGmNAcBu22GTE3aTJh5wxgnTA+oIiiD7wA/kwukZKA30V8YXc
QqLNEYH9Erw9hxo9IM2xrHvUTth5OFqVw3Ls6qul1gRZMOgbdH/25zQYCG/yDtGT
/KC+kDJHkSy5LV2GHUWfsRVBCDCZs/7pClu/XECgbjhyaV9enNS8mSwji8Nxy+3u
ad7ZL3ai7brs5xXvpIlTuwOggtLlAXd76tmMbgdV06WvV0A2vyh9uEgUG0dXfoBU
But7jsc7Qhj2wl/GyBIdxeoz3T3It+v0n0ApyEvHbLs8EqahgyPh6llvKJ2FOtTJ
mvPro8wCXlxi54tvfMx7OqYvtDgZ79WBCPodKcm8NtS4yGWKR/aQDCcHKy4CefmW
2ec1I1RGpf5PpfiFO33p35gRpQ5pYAUdwgL6EFhkwoy/PHuvZkD5iBPEVzTzl4oK
QyKuq591k/xZxhGaXbWRX+1rxPpGiGEpxLXlHiocC8X6fzHKXz3ZSq2a9TCc0kZi
6LWj70gFL08n9u46Sf/K3ZjQszqBP2kAfhQSZqaECSU9lftgbWXnKuabY2ClMPsR
ZOXP5PsUQSNfXV0Ovix0Cnujzuk9Ph2uAI9o2yBBseotXrspZY9KZTJGXlDMtgig
0eHgMYSfkiPX/hFTECa93jsWg7P3mpDhBvGhm/SEBTrVFqAB+nYVzgHcYy0OfnOs
jLrEncYZiJvDie2fHPlyfrZVrZPRUp1+VUckkcaIajQQFu98g9TCG1FFao92yR2d
kJ0xjARh1bjImR5AHFtH0q5Nmfa2Gb4jr0D7eL3+kbbYxTyHK971pxtQDJGDN8Aw
LjM/WkQ4rb2XA+QQjIzJxw7aM++WU9OEKYSr9yh3o0ESj7gSnpJJolEPeqQNCHmL
YuW0KEtA2FfywZ89AQsXubDtH2d9NSwh503JxdeBMWVzeCsqSYD0K33dyTR7eMiq
Z8rCaBbklLGzob4rp2t7/Jk9FV9iCX853IafA+suJLlmYJBy8vWe1VnvDax95tc1
ej2+72JLhUiBlGbGzAusD5z2xCjfZGpjQcb2Vj+H/PDkwDoUNzvE025yLGMB0/g3
SV2+3FXB3JfODNoeuZtsQYefpZtTbR6XtIBArLR6HqEh7t2TcqJIfBuWR0IGInTX
sMGEXnoiUtkvH2n5GflQcNl4G6kwVS8JAdG3xa3gmGzeopJeaJg5YKG2QaD7XkPy
pH/Rj8UDCuV07ZUXR4Nv13DE2rX8vispBaUg1d/Z6SyCMxBqe8UrljEJLr6D9wV2
mCs/A8BKvDeGjisSpPglnJeMwH3C0NRB9R6557Pvd7VMa4OcNdBqMdkw/ExrUVTT
WyfD47umg9vjK6jhmu6K5h4WRl2i7lecihdLcUWBa3zSzpHNRDQRieXcpYCl1q83
K7o5zl0n4ufqyukhG/W6KiENr3dVitOMJUeOI6ho2ZAkhYgwkx3PcBegmeDARRLN
kjVIRWqq2/axC05K07aLA/1cjiCPVAWatZSq3y/Fe/0qLkmjt7wrytK3LzNQPpzn
wyYlQDzoOBaExte/xHxMBwLZAPMitc+GSHXsqjRR5bYzgblp9ycGROHB2jk+F79G
JDUJZZybuvZascje/9hnpqNUADWt/gy6nOjkPApe9oS3gJ13jiBjYtmVvSJhQBDh
niPXiYtr4uKSwzvp6HJ4A8Im9yl103QRH4XbA4WNtH0ZE7jXn0Nucq5NR/wTShnR
iT2bBiYZBLP7E1qVFlwTNE4t6l9AGFsXqGthk1aVe3iCWZO1NL84QiTpWyjtd0pg
vza4wetORuOKHXUyFlnpnKje/JK2dDpx9H8bAL/h7sMfiqGmJPArZE0EZBZiV1Kn
TcjDqYEWqBZCzIa/4QpMiKFscIcmH4lEL8Oe49x8ciucQf2qNgdC73DGsGKy9N6x
AJflx/MFACCXFv6ub2w3c7oNoOgWw9L8FfIEEKg29iQIPwN42rwdi/pHqtzIW1Kz
lbXrtXUppbZlC5Zf7TYQAVXSvDrF+ZumPojfVpzkyMYgpj53ut4cF8AId8wPxGVv
R75QosPC/GHiX7AdTWe1A7TTJ0AULqIno39LO7CdhLMy1BGVFGI1GKws1z5byh/U
9MgDVImJprcbNkNUCPWNdNCP5BE4JHjXCpjbC/GrFIGwSSoraoBxHJwUsKaoeXHe
tpSJ35lgHPo9/6lPwudTOPuVmocHEsdqOEwXC2fFUSMei40BBSZPd9+pNUd0t3ou
stsD1sekL9rqMAmvFgQBet7fyPRbANxnjS6Ibjb12/3sfuib/wpFGgkaEPV9fvwX
v/wdVQxeqqxfm+K7i73Y4RGnjUQ4FoiaoS2vAUIJDJQA6hQoXoJh97MM1Nd7M4Es
w+pQugdpTmwAnKNnjz1ggBOJ8TDhy8LNa0lK/b9cUP3OwTV9FVIFVOzcf3kizKNq
PMiG8NO5178Olb5AIkRJjfXj1vi5w7AVMFNwwGXQHHYpXP5PJFGHwZ8H9L9FwW2s
3d/lr7bpdFJXMNCn94Gj8zZZCeQsBfuD5xulZQ+3M5CRG08XvGqueTsMZ+vCZ8Hw
pgM3cw0tfEHQ5ZOGX6klZZX5L09Hhnq2poUMJLKCE9MhAnDLjowkGR+HA1ykYY2e
wn3OsqJaAV4bqXtRhEEeWzlqjSrIqIClwZzbxqvWUiaBSUy6GFHvBnHRf43UKcvN
ZVMFB+8Rezd/Dpv5bEmXyyEJiTXdncdfBw/NwGJh56MFOPoh2TCRJDB3mJZsq9bF
MZzqeUR1ivHerYeQbrYlgUYP1AEUhBOpNKNjScvfpd8tVSwsMHtZ5518mCLtzv5T
9nm2TrDaw5PMnby75QjaZ+pQ7UrPY4PKHJz5gLi81Xk5Ztwot/PFvWFcsKV1rP2+
arPLXYa2n4wqlKcggOnVo2hc54SPwB90sGJGYgWNKfuy502ZuFoCjMpB7x1JBIzG
+rb6Q/UxtZm5ihoEq2bXm1HHUF1DVeZSYG97QohPTrg/DjS3MHjgqTh1IiSE0Ikw
noVG/XlXxQBzv+qJV7HtFlMc+lxqhCvqpdbgNCNn9vJqNhiz6LExtWZSqF4iHDsO
RKzMRgInAWlFj+dYB2/xotwGWf5PIYIrp/B7urAnNnicvOUSkuAcHvlAVd5LiSyC
G2bQ9QAi1zvqMFtABjZe2EHI51Vgy8+mx3mDprP36ULnEkmSqis18Zvgl91EUOEa
pI2y28JSohuO1NG+shBUvh4P4C/6RtJ5idcOIaih2BoiDc3cHs72FQ5C5R0Iu6v6
MVhMOVlcBiX2bhjB/hEHJs+qzBcEuicAkPGUga9rGpvsac10NXVGfULm2abW0TOh
QawKVi92uBZgMlzhlDoK/vY0ouJpHmpw97mlRybwM41q2GDoSvZPYdBSOewrFeOp
VxlbRF5IW0g1cbSTpjLQZYTx0PbamkowQDPB8Nf9IVe2LO+eGnYe/JT8l4zVRFTD
eoeCfUMnCwkojrk9zTOE7PEw4+DdyyUAE4vLBTYQwqndka1hlqoO+bHy/QtYd/bw
Wd2sZ2RZL/BqCW6whRmLLSNI327iXFJZ98VxuskLglgfkQzOdkiSzLdaiE6AIbFn
yR0x9oP+YO/8zQnaEHOqro7c0VGtCEeH3Af9CbZuceWuprF5WzBxa0f19aFmdViN
YqcjSll2p0/ivdBwWCIGfo408TphO+qZs/hgC61qcHKTxfig0OvCyH7PNllFMHbU
3yZv2MV3YO8i6MhzFr/BypPHEzfkOctFVPrK2M4df6SrHpd/UYXqvuFiIu62Pf90
rnOE/xVWlfRBFZl15g1F1yxvcN7F5EO8bIvd6ZdnWQYq1owqvynzUfjJUCNqDp9K
qt7rBdMGah80MX1zeD8zcbbQQcimeE09MJTEvOL3vnhE3wbEmOTGBLVOW/osi5/D
7YZ9XZv9VB7L4vdQOOZaZ7VYxbPDtVvh0PumQkFPE5k84IF0hU+7xy1AqiI1RcXG
xwPCUyMTwSNL9mEOEJQWzZcX0dWFlEiNQFL9jiRObrr2a4F5yLdCYUsGVprjUZFg
Y66Zr+7URCiaVtVI5rqO4d3G0rcnE9/aNCBhxTkMWvLOh1nvT+a+nGBipOWF9Gme
RKQgNczgiZV6Bxzv52mitRHJ5EfrLZ3DpTKMj6CsD52wSBWgeAgASYFW/e9BPlbG
w57uIV6Mnzxm0UZpIdLvZaHgaVd8/8Ra59Qc13yhhWCx58OxHzBM41ecuAhOJCYg
b03cF6aECRHw7nDID8F/zBRyH3h0lxSXCDJOVjZZMIjK4EZMZkNcSB+7w5yN9NU/
Zpbzlx8XCYJb7iuwScsQYn9DpzOVIRiPZdKPaC27RT1m4HfitfvMmRqeyMYJIlTX
cOk2NKs6Xj3JYgRkSlpR/VvBmRx3rRnCHPPMoMMqfv+1PdyXQsKhnRwcB2/vy2Wr
f3dy5ug05FU97zb0nNpXZmV042XIKB3DItpFzepRIXxr0Mx8Ct8ep14s09WMD8P8
dCnurItvW2FNZhdhe16hDcG4NtXrBhVlZlEVhabnbUO/VRbliq4Uzldjf+b2WTQX
OZul06N83TKOxwMtAec1/Qf5JpTGjcQbv1tRoQwoqM3RWVAc8pc5+zfkZkX80YIB
wTSYUdGWzM7JV5rH39Fi6fzSY+97mPkXPOA8jlKSSLyfmEYBQj0u9CGYywFuZH7G
tFUTzxeu2b9wpVI+zTU4UVhWlJfkvbhHAvUu8u9EMECg/3tH8i6mFOg1FmGiwZtD
BEjTzgy9W07RjEVQkZtng72SL9H1s0J82DcY9/2Z9Ina7gziPjY2OJnd97mxka0j
xy8pT6jVt6l6v0PlIejTx14VK9BJggLOMVm64hReh4TWCqUMgu2ZoFrLih11NgXh
O6z3JdNAjm6ROqGTzcAdlek/NJZLYPETBI4I7CE/KSAWoePyMiLBn1tlWnfMLegb
1cOYBZDMdBPSCsA+yZSFh6UUXZrcpxrxMSpKZOftZJq5SuyLmCN9OmTz2mIYnjfy
Qt7To39ogw2+AboJnJ9avW7CIRZI9j7+3JNVv+Y00CgSSZZec9UOAaClZjC37DDt
lIAtUiCk8dUryqIQKNWaSkdfOKzt2MIWhAf0nwVm6LCCMyX3l0M5XepksIEp6Epq
nAKS3iOytq6vhwMzzKwpmfGJdulnPSfQ7LUC46iD0j1x7qkWUwEvmcRa0PlnPhuC
4egqAI7OwJmc/l5ZatQBWh5O1MCusv489aAnrgkHB1Wcj7mlJecs23h7S5uf7PT9
LIaW8eac007VCDIn/4gvM4BOuYWweM2QbZoEjSEYM7FzVaz2oDPvxjqSlcQaNg4r
s2GxrpLOgFYByfrXQctYiW9d9fRD0Vy1mhy9O5FMT0OPYP5/LaFPkJhzQniNTo1A
16O3VmRe7x7ff3gXIA2oIJfTSXaNsA77WDh2l3EKyA/DI1mSl5gqDMWS+/XTI1fi
a5TUBDlkasAFI/uutds32kX/tj6zO9D0nN2Wcz3guM6qfK1EHE6B+9FhEWi/dEHV
u277G1w1O+r+E/hqGg6PC4V/ibuAA87AvBW/lGislTApzdKivxSygNG2AZMZ0WtI
hBRvblxQpTe0o7s798nkShlHhBN9sPSwhhgutCc27R15IZOKiAftsCJJ4oAvvU7A
CGtLa78o+QpX0MWJvayS/GjqEPEr8xsN6mlMDW9Djrer5lFxp+rTjcb7ZAFxlyC2
wwfeaspivNDo6ua4o0v/sMaJ5JlGir8pOV52tR5qaGKtcMSwsYZeWJwjDo6gOPVt
k1yjSN0il2z/FgjTN8GTdqVocMZWkT5zSqSVX1I50mYbLuoozFAqE43I5P25UrFT
m665wIZ4yjOFepyPg7AboV8zML7Z0OxXAv+c394v66r71BJkm9lvCkU0FDogM+FN
sAAeHfMGyEJeIVgjyLcbHVHRqoaXM2czGFkrYn5GeBpxOWDz/T7ERjMZm6QNskt1
LFhDPc/GL/Ggjb6PYZv57oNcRky0fcPcV+W9GPfkLZ1Dx595JZxOawbEIQzgdmds
g3VbjcxUafLm7o8YHnsaVNGSqx3tIRFFoHj6dz8qCvKO/LrXPF3JKOrLKI7QylJP
JEgKPEeHdMlWMYdhCOzZftTTcK6vd0de8Ej7ToK9+saeBibcYIJDvdmWXGtCD/W8
eGRzDtCKWjiwe01THKv2oV2z/jryyXwgJLphhQofi+srRJHnt0SRm/sQQbzQuVsQ
um1d94P4UPDjeXgcHAfJo01lwhag42TuEVDuOZ0Hfc8131wfNxwlOIBPo/kpm6k8
x0FNQfkveaBIcmmhibQjJ4FkDmKxQTbufIXBPNwiZU7Gz/45h0PHayFNynLZxdpK
PbTopCaviRGjGqFF4Pp/9bY1Gr7suihZTMFtSR+ten9B7nC/a0yTMEGtF6HhXW5U
h2mivA7RB9nHSoKSR9RycdtEWMjoY6zAj63nXVyFNOSx3bcSUtiLMiSw468+ig1L
Q+kEi8NrNn3bnjBhca5O8uhTYNI8QWA3vhq3BqpmPVLt3MKQ8mayVZFfjnkgb8fw
PhXNjTbQqnVZqEzvWMPhiMtDKA6TXJVf6COUjdZ0EpD+Sx+LRyJhZK3XpliTONbH
/U/FnkdHVd65i3aeGTZGSLLKWSXP85GNcKmLoXJyslagrcnDcTopwZmYaJUscY7h
u/F2BkOU7m/o12KMRFe5v1N/J2YyEpEWwDvJWItQldahxtFovk+Lrtl8GJ/8RCj3
sUIUhawDVlVvl5rzDIakyHvqHlFKQOFDRFw2MUNnzlnJgRdymK7SoRy+CUopZSkt
MUEqt47r/2q0myBLOkTSNrV265JSOKqbUvtPUdWAGp25mP99YdvnzvNKhNHfNt6Z
uMjya2nIX9qu6mY7CqNEmWEv69N8CRUl96Q2R/iP5QP8hF4B6EqFoGrB1Q1QHkFa
l4/je3O9ydq9/nvDIhNxfZIgjMZbKcNiyDVlz244AorYxIon1oQx/X6OrIGTsdDL
t9BGU+WDpKN/n2Cgx6VQZDSmSNpO9P+4MZXMJtLrunyq6loOeAvq+SZjteJ5SfZ0
i9m2pq60oKKPR3cId+uUUYeseyVdp6ylyno//6mWSo6LESewNVIVbq3YJSaQ7rol
AnUhzVHz49+1iXBlWQxxGwrAdKWDkPnl7fab+LdGjSKkW7MehT8yP1jYs3rR0Dys
S+mBwG7lIdngk9u32IVO8nSqgCqDEw5WO3vD8UuOl3DrlDXsCbzurmEOWtNSiRMw
MpFYUiBEV+2Jjn3HH12S76c0D3eGoiyOK3r/Ia/INmPhgzJNl5gtYn++gJFRcEyv
wAoEvV0AcLlQGhcvMQQJ6f/gcUSVxMxyuD3pmgQJdO/JuLGjq8jS5A+yghfWJyrm
nd4YEprgoB/vOuVsQ8gcr6uA4ihQF/H+2VRjuCrC1uSPTd+wA46IBa2UKuqU6vLr
+OLk5thZcyoh8bjbeln0P/qq59cgxoUNjW1JUTk1BHRGvad/8BkKctP0qyUl5FcX
KO6jxOrrEGmTT4xsTxxPkNRoz7G0/Du117r4cBW7yc7Ckq26Ob7rrBS/azsTWKAC
5aCGxOIhVVldH5iB3+CgZoIZCaPiKBUZDlXWuX6ImsbzqJjNb9iUFdE2rUlyVEj4
nIOP75GqZCEN70pSNvQ3DyYaSwqzN/I/oNs5DjkSmOfa5RZgiGQ00CRSpiFc1bbg
6YAeSdQQWMokNRBwNwS+FDqoFYcjBUqOhVtN53fAmxiRW2TXLXLVj6dWzsjqRp62
dYRiuuaEy6f6g/4WjiZ55zBVXfCOvvvausD5na9fSdcnKsDX12dOPwXjLvYX8rwM
yC8IkLDVm5hbg1Z83LiB0ImkDVr4zrRyomutPeONk7NKVaXi06pu7YR81kFVVQM1
JeSOdtTCTRL0BSanyZFJ6ttCUQf9k8u/wJkkP0gJFyuK4B6IIbe9Ua/atptEMY+w
aLDa+uVvvEdtO+4YBNOEmbxrzTzKuflydIq3uvGH5s/cIJgEspvzMIr4S4qs+cuH
6iKIPgPlJRns7WKmfqQmSFhwreaAc0ZHx/9ZCW3CgdW55rQ5CYw7pXrQpobBmzbh
tPSoTquIBee+TjiaVe/IryVc0nXW17XUqb7Ycwp1z5Aa8K8fDQl4Ji1XD8vADXB2
phr+5/6Afzgn/fGBANyF+nl78xwGoBvQ1ksIHpVE5tikTWFE8RZCZpqAqliuCX1S
YoS/No4h8UHOPeEyVWYoEHPF2/rg0tTTUw2viGCtlYiQ/YS69SrtWnvgkoCGzBsO
kWOTorGWM+m+lhrxKKKjOI/vLZcCPNF7ZcTWMxFIj9Wdihfk0jg+j4uaO1H9puCN
tUnMEdnuu8ak1rMVsQ9xz5WzlOTsxskbWnqlUHTZEdRdMzxO0zKWKXKiOZnwXypE
/GBhr2L9k6L2WwPf41P26ngrAIYTp+bkRKAn0RpcxznLg6ORN18NvE6WNV0mp0dB
ex0FS5W8B8UB0uJ4p8OReImLWTOnRWCsB2wgql/Ws+gt9I3QiKrIKyojf9mCytjR
8ZM/4D8U6cep55nJ/ePuxElZBOs+frc91kz8Wp3yIlA/csIC2Y1zVb6XtCqCZSmj
ick6EYN/TkTnimH2nBdVMk2KiNXprF/5LT4odJeG+4XPQBxlCcDAEsdmKYx7zRv2
ZBIznZ+dnxGSl/pLcXBEt1Col4JGfHUC/VDPL3mXzrQGOh16UK0xB/CthbJNDuIV
IQQh3Hph/t6tZv0dVlpKv3HnsiCwxZBi+ruyTCtNhabrH4M/y+GeGtp6QrYcy4fu
KkbpD0YRc1fmnik6D3P6shCLs6k/uaOVfDRzLKrBaUCvMncaaWBJGJSWNAe71VBU
cAgAo2SuF4GOCDl9Qzkl3dcPuFrrlj9ULe80lvtWQhCrdpNMWmOMafZg2p58MXXA
BE3vyLfi9fP5btKoA6HtqOTWMpSjW0n8uCsj3EKIxkBjpEeRyY6vyyTM7stCEBJz
8wmy8g++nB4naLm3FzxyigG/bI16+xQnZCdgxsyoSthAlM512tG0lxsgok2Hb9qY
a2unx6eXMKfv8eJT3me2unjVhRiXa7sjlnaW7R9mLdyCOy7LXIUVaIv2lEIKsk95
V80s95w0YuGalQpamv4udLbZcHHk4Zst9aPIoJ4eaprEQSL2kJXgteJ/eK9RE5VA
W7dV9hsBuAr1PL3LdLNSBKknsnZvKyGZODEIggK6TXrZWwAQfwrioGQF6HMJKM1T
2Wv6xJdaDZmHZi9ZZEU4xvylUk7r4pcpg5Wuw7dZiQCo2zBpAyYsqKSLQpwAK/F/
R4Ly5SpCud4sfKcHoL4YAr+vcYoBg1UmPiywWIkUh+htYO4qDCXgGn49RjGcBswF
8J+5DFJh+hhT8xOJGYJKevn8Ldvsv6eNCLHAbrk8ejJvx5cqlkNv/MTXXHdWFYjI
YYuyFhRXypg9T6U+MSvd3VHtpRIToGYLRlSslexOcORRBy6OP0SvX3nhAsb7b53L
z2BMKyZHVCfAUZWJ3H4AENsJZaimmmqgXUbcdnwFHb4oUxRQw+vND8Lvsgbb26C4
8v+UDspskj+hAar/sLHi+EHh7PJmwbIbu9b4NkTV55QhqNq4Y5AxuS3YYGTkRyKL
J5/VNDzX+2xPx7h9p5fkOuVj9c8UMUfTYrbze+3GXyDkPwwFFEHAxdi7vnQQQQ21
+4rRa24SMHd5whhXH/TpRGQQwnVWM42anuJY3bVD9G4meSNzqBIdxQRHzxeBeVjX
2SkE7uaj4RROZzpqMDRZkF2adwa1+wCsM7kDiFJfp0Z/j5l3X2XiGVZYBt6fr+ac
cj3bxZMc1V6WNiRszwWUig7/mt1RbndVRFOmS59zypYybRHdT24meCzjameJc4X9
o+WbUCsCh0n4ZpbE22TVDXfUTnMUTN3ZONUdO7zQOnwFB99Obb30K9bB1ieoOwUO
p6xmUjLNNb2JwCFrV2yu0BgXDswMJGlFbjOHaCguhopy3QNUlZRYT968cJY6RE6W
qqRLhL96dvzz3yCwArQoyHfV6whkGYSxm/NMn5sd8HoXXsTndnfTytKykApVdJFH
jj3ovtRA2gA42Wf7d0wbBOc/BdT9uUBJ5h5zzs2V9R8Y7BbH3p/AN1h+TYaSbC6r
Qa2xBL26hJ1/dWm6sBpG13ivT9OKwRjpWdTUVBR8gAUak3lVK9JSfkwlAcAWqD4Z
zDLgsv8EcLA3vXVH4RrtR4D2GBXIthiiz748XqUwLIwF/BJA+LBMvZb81rBQ/+qp
uuQmfeneAsyPkeWTIweb8kKn4/lZToB9YkCQAYxhPW5UIGYvqi5lAQ0K0fF0x5Dh
W9enheLcupRrlkTLonnHJmwvm4+LHouDNSL7N3BQKaLb/wBxNySt4QMkbEq9uPtM
QiOEAXBJp4gxVspJTEVwgFsghaLO+UdlEbgMLMDV7vGuHaxrIxe5taWZu4Z0CNYd
roZLm6+J0w9S4OtFFKGfuUzklqCeb/IwG/NTryCkEKXLYb41lT7s2HgB/rpA7nqk
9Kkw8XXzpA76NlaEBvHvX94y1wJBzDZ9/wsnQsbJZznPm3gLkhlT+yqh5EJ7r8pI
SKWTmR2VRsoZcWKMDv8UReWf295bXMHZH47AxR5gV/XYIIdjJ6Vj7a2unfz1Bqr3
NhGAzIBq1N1FS472RGlyp0GwsvJSFVIseLLZ/RK7ZLCTH84US4lSQDqCQmvELJiF
rv8ftkVe3QGI7rh7NX4zyd0FqrRA5/1LFmWPHH1vgdPoVpHcCRVpcN+q7rCtDLGj
y1IHGgOPIUywAJESnYHEhmEyaoSkSzCh4QrSaeDKMPp4ephpd+DLv4RFSP3pF+Qf
NHor6bZ6lK25tdMvuw8qzDKM1/11eh1fK7gnSY3ti9jfvtqtbe3Nyg0T68UVC34h
hfeOpoV5gDk/ZuKrNoY+O3697cdQQWgyiLx9+T4YWlPFsSAFggcMMsXDQJIKpuJ8
IiRIUSHYxxluwAaEizwbgcYk+45TTkRvX8dXaGnO0HHJ9cN4pqXvT8qbXWNqG559
nyAZaZZChA95xcDKNS31cRxx2tEoFOyQLW5WysKv+kjPtCgg9bAoKwR2H0xIIV7s
bVwNAg9LVDQZPwtl4rA/Ldid8I5jvaG+Gls7dYfDwez+Vb9uduUYAl3Ub3+hzhIz
G+tFDKKJa9yKcQPRNJWMJyRl166ew0yV+Ah/kBR6fttyK4pUH1TrVK1VPRRe+bTB
Irl1qJo43z+KUC128vLSmSEw80raHwe4KT2csee+SCHWAojgC5WCtUhkT2shV+Sy
oUEVMdg0cL2gfMqSwi6Gn7T0gmk6a8MYt7Y+wCMub1V69aDM5zj4Gcfe4lGlQVys
ql5Ikfuj/usXfeTtcS9W9OU/un1vt+VKNdRLFIjS8n9BCB9kUTbY+CxXBrBSkO0K
PuNK6Qa4OibssKwhStDLp3wA9YUX2eYKoaZ2L27PvktvZWxpvmctvy76YRXlC/mT
B9hhN89VKBXZ+4cqo2sLRL1KaPPOxS76xfYQ4gy6tQNPTA6z/5cKlgByfFzI9b2h
uxoMz/26f9Op0N+RfrqdjZgdCZHce9rDwWEsUnUUIya5a9YqF8iXBYyN9b9dIUnY
6jfgwDU4rFMdVZMxhGaCvnIQKgo8ppph29t0oSZhPYnpvvohOkdTFpg/lVnKKGmH
RkKROU7cR1TAl5eKNZ3XQXzUINBFfcv9+Du0tR2LKrIoFBHV6Z+Km8kBpMzw/06q
NU0DwmXKv3mAPHnJEBmF7DR2zZU4YT3jI1y4zML6X6kDkbsLfGWeryX6bC6bTcyo
EcxMHY4AOWfYY3bIEh26IOURcoOadDk0STcd9VR4fIdovA6FdlE6L1uPR2wi99qj
Nbz7hS0M0Nlp00wj450nnOdp1LAlxD8ovNSWWAMIUJMJP/rWKGm0M28h5lrdM+NQ
75boHlqZD9RL6bbwgkk5TpcTjdxALwYZTncvuBy8IADuFAKA8XVoAU9euZVCUm2J
YqEh0Dx/8qDS7ZrQwEnDj2C3ByqmfUxAYUAYoRu+Ibb142NgedVk+n51VrermB3L
agw+jjGELtDbg8oymldGlBY/GA/XYY2R8mPLbFSTJHvYe56zyI23ZV6AKD1C9TAO
wSlG470+y0VZb8+HIANbHkty8/9rpQRBKVJ/fcUvoa2my4HgB/GbVMRbkjToADtS
HCtg7TNByvfQPso2sSq0Q7pgRFkyFr5DjDRTChKq0c1bMnQbaIjJUjdKcPEs5LJC
ClN3p3UzC1YC1N+4SnTDBXEArPesiBXcjd4up5qKh5rfH47Ky6kcmS7U5x7GA8Cu
34Keh8lBrXR6CK0cG9/r44nUh9X5mU12UIWmyTXIXvzIicIrfnz2mqCiD9UtWNM5
04gm1lGttbLiVW1OQB+VzKEQ6NfFDEtZ2/xYHdZu6sPG8SCiIaLvIlXAO2fSu0UJ
53te3dIqy9VjmexmtQSHvpeBhnL0y0V01KrX7m3WF+Tb3CuqrF/gxGCQKEn2kfio
JX11OfBklptVY+iI8CFlWVfSOiVCtp0A34HgnIqGc1OQnx+xoHfVqXJWNp2P1m1u
nKZb9K4FRPK/PFYneB8W7FUEdUkIKr18TNXx+kSL95DwBGBy/UapkUyhAObmTwHy
2KPc6ktiVuumehlgqsRuJ7BpOvKkNkYeHoCiUC2dOpACkk7y34S22Q7viUUKSdXr
XRztYBt0bs/nkL/c3SZ4uO1Pq7EFJ0U5F9kC/4SaMDrsIvgdr/EndZVZvDJA0Qj4
IrYECYoqh6derqKnV4xXi+JKO/b5mOpTTJbufOUtfsk5/0KJ1+PzVAopXQxtF1n7
IwQyBly4ialj3mkGHKuQ7o1xvBB97vmF78EbZGf81luaLtqdQcsFHjw2DaNkyIcv
eXuxzBRSTLvtTDx3x+6QTOkNaNX9my+l12xkl6zwawO6nmFlUkLiwv34cPAXWown
AcmSzw45epqNR0Kcth0/kx1aEAfT5AztZx7IjZYtR6hx0QzTNta+9fX2fReaEQad
zqvBiCJ4RMig02BLFDFPhrx/O81SzNg1/fyTEzi1MBkjEGO+Zf2dJQQJJ33zG95I
qqC5Gl9PSqOmOo2jm3dk/5oUGyiCYChK2SsAgBFtIzNCWrkhkqu2u44dpBF7CEhi
2yh3y8usOpJwfHJpbsr7w2emVjj+9I96IWh0mOQf7o1e7zVu+ePDdO6V/i/PvjiY
XP18EelrIjmduXF/1wu17jUYmbYoLCGN6Njqv8C73ODZuOcfYsDjpfpSrMx8d1uM
0bU1fK/bts40DzBMAV8sgsIK6T3WEjf8VrlbRXcVcymDJIFtrMhjJMoT+qgNVlRr
OC3krsR18tAZfujHthiAXaX0Vh4TsbcnrfoIXcPpWb+tn3G9BMWg+5D6XwQwCUrP
OACUJN0hABcrBar6R05qxj7nq0gKPNgDK7WXHoWrGnO6bx+0hR72l1OSiaSxXAQB
WAjxIPag2821GZnhpAJ7f75Zj6NKBNt+AqzWQZR70u1/MNDn1XCB9f2F3Qyqp1MT
UpPl8SBi3uQ/mpIkLt8v5//FIGo+lN7ASFjI31eV+UIY0orQDfHPDyP1oX9bbx2u
9nkBHW2tL+tBT16D4qqR4vOwGBSBk5u4QXz4TUAIAXdFWwbdCbLhk9R3CvAlu5UT
Cxsjn2tFPV2bHOLDeXVOeyW2M8z/1zweGJVob8zb7QENhCDSC0M3h+KCiPcr3/HE
+dxsSulhgdqs493khk5NK1mvXS/Iqvvkd/ltaMFPWwLAugDxtXLTYwQkBLgi6jBL
SC1+IJG5rIZQst24GnIhZMivi2iHWVRUAEDw4qQG7T0LYJYTZADHd5enWF8maxGd
PfI/oPe2p3ODoLArIlsaHEtSOF/hLrcOFc2GZPlp0aFtbM9g4vYD1p6/xNDC/BuV
tvFqh0R968lYLFjSW7R2IO5LAmQ2zNa6Jv0TKVLvDqoToN8uo6z4H1cB1mzlfkQ/
Fk1gqQdrf8nuUdoQ5bzeWDTiZaQ8JTQ8OzHRC1oSoP9v8wQDwH04+KiM84a3FVKS
Nc6IZrDCtbRk9tO1CnysKpTfjvaymnsTF4zwzIGnRPviympcUyCobGfY9fhoS8wN
CRXhMD8n7UkFxLU7cPHPw7w2OKLQXYYf0EWTpysavwOvuYhNB2WJ0ostLL+cUEK4
q3AJeamMEnb6XGbFWhRsNV27sdzZiLOJA5/I7iHc4VexldpgY67gkE81Nz98+KGZ
KXR9MkcI8yDi1cRkU9CMWneMVS7WgY6kDJVu4OI4vEneU29L1iKhn0wXJVeRNj4W
E5dEkiSYkKAkhqBcz5mDW+0gr1sVULaxeagp0WaXFz/3lBhVdr0OcCp/fFLqpSGC
shG4brvJqtG5jJvpt1VE7RhUXuaTRKv2cIdI+WwMB3zyOO6RafARV7+UZDtrcS9b
9otmFwY4TkcqLLnH+xwzEuYxu9d6Iq62nUr5p2QrLC/L6cqogkz9GFAI+o0eTPds
2uq410sSX0FIpDnrpNQGTjL4WynGNHwJ7ehxiCJOhMdUxbTnVU0tQGEYecN8oQKK
PMmOBYKFJjmPmpYpLVhW9IatAZPhbPL1CKWAoCZoaSpZVilQpCa2jh6lhRvtoGbM
aeJgg3LtfWQZGaXt9AsXghSsoX6bcoqH5+nUxWz7Cm3g/PWHIOuxP6rkl9E95EB0
QjCUcPEtWyMhosrJLOEEPo0VwkYf/kfynvfCVz7DRPBskPmz795V6R0+Ou51Scdt
a6ZBX2RVWQr9O5y3hA2h/HIieCD7/G4kHoLn4QbJ3JCVLzwNV7gAby6u7mSV8gA6
8YwvFvOyXq+6CwLDpAL+/afIcmw7IYoRHwY8aWHY77nABjF4zkNEwIQagXPmZKjw
/L41on8wNkg5CUuDq+aDsmkFT02Ff550r9KuUIT6hRSbP6jZ5bfwOVdCaZDkk9TJ
0hBEi0TSOCAKAxuw1re0yXW5mbQQMA316laeiOUk1FMOoQhd+IoYOIGLYf4ZjGit
MHaTcUnfhVmHXoNrnTAFkBbqiixqE7pJxmltBlP/ERgfThJYQN5FF0GBbpSlTdix
pOZPL1i1HvwV64Uj4qbIzM5fYvDhV1a7XliQ8kv3+u1nHs9XOTLD2MqcRd9DD2G+
zRMEgp8dfAa04C9MY5kUuZ3V1dng599Oy++X0E7e1Znp+tvLOhD4Zm57LuE8zSfq
mRQH60Xlbsd+ofscYs3jQyuH3um3KpEEBYS/wPpbHexQJGiXKfLWzcqYnIjFBky3
Ekd6TsC0RG3pcFR104JUOSGZ5s0lCl+jdu6+U642+GG2JsvpRobfdYqktK/5bTbN
MQYW9clWAUxM38yuohWHkg5/1gTcGdk9wr9SbSHdM9aGYb2FdA91lxjK3fhhahDW
JyPfFZ0kY2MvEa1lAV6+nq8gqc1xK0zZcvvLCRRKZiyzWlehIfR2VoSsHF6CBULD
k+zr7P88GspbQ+8Z4IX3KaDOnqyCNYbQX8J4aT/cxPJPNkmjIRmcX89jhJ4qQzfl
Ma9LjYMZ/EuIOo9VewXem8EZpml0nnJzszyS+zab9SMqIbdUz20upr42Du/GdKM0
JfPUtGEJFNfJpDpkikgXAMP5U3Gt9K1xBKB3mGnYcS/3Y/k3w/7EQ8C/XJ/CTzQs
gpnbvcSNwJx654Mc2BWt/Y/Twusj8GqWkjFNS5JQTpJY0bpR7eMXxavftKvMnJQr
YOJgbMDvn07evZp1dcxPadBexB+W8ekb4BbllJOBxwU4GwwIxQ8sg1DkEOFKit6e
Z8z8hgSJEOkHwbZ7/QaPjRHdPj7iPLJhx//vEtF4SDbr8sV5r7QFFSHbpVB+QmGH
Ac8SJqYWAOZ8tqS8rfpy/q7ytQliFZpzNNurlxSgFidylfdUoTJpitd5bDapDx3w
a99maGDQyZZoCbwWHsBp012fkzfW61L3vpm2vP7tFmrdIJzaI7AQYD7oTDiC8ktC
wNbRnhRjVCSgnM2ZQEpHBIGvfcvq4y4qip4N+YXjdCMzkVXhViHrFUxA1OkmeokY
d/EWn7FyZ4yeQFVdFyQZx9dzYVJSgzHZtR+q82LL+o+HT8y4Xja5y7VcpzQoQ3RF
OCcO0ciij7DCB9e/vqN8llI4PQuJKM2npS2uElRtsruD2H/RH2kRMwit5WxOv7h/
E8jNIjK85HXZ/asL8TslEAJOwmdqXQD3BiFYIwi9cViieMrMWGWzDbU6ccGjn77T
RaKmXZBCFVI5NDiIXXM5JD5Z/GtEWs4RbZEU4rY2prb//gTxGUoQkCnLfLpRVoi3
PrIdwykBvN3u/RNNsVW7aR+luHTGanppQm/Fzsf6lPlzIvO+oaBy1rv/7xHo5iiq
IotLGoceGjeQilMLtoqlFsVRnHiRYoYzGE7qOfJc636jeknCgz/N/091NzPmpS4V
5FRNNhyr55v0ctdSKYq/+Zf5HsteSlC1j6/uOEYJBTSGcBhk99m2s9pbl+hKUqsK
blYsBYAZEgBRVjvJuxTRwhtVignDOtOiLN+AZ1d9a7fM0NCMrc3+1NP5nNSnSfhS
qpqE8OMq2fxC8rWbBZ6RhAaLOIotP3ty7C9klgIFK16NfLYOOGOQB9o5VqNy97el
8Nm6Yoay4YvMZTBEvGqQCSDndzaJ/PeOv39PFXxSQad/WNBwjcAz7EYcwtG0m0qy
H9rx3/8C00CW8+5eDLdL6c/PiI2SV+CPssQsgjTQ/q4L8UYp1uHND1lqmVe7jy2q
fid0dsWDpwMaml9svF66vKoj7CVweypIBCDgG2fkHTSdUc7xep7cqal8KOBPQjl9
p+yY5fxeVMNLX5dOjqHmQxFiouWu4Nqgx0e2FwxQOuc3OYNgX+oMYLItUWFtZlD1
4v3Tjr2DWvEzTrlni7JYuXYipdEkz9Kssyzbwat6jp3bQT3+0xiNRMkXGAbOx7BO
Te0p6fOrWy7up3SumjTTq+q2TbHYWbXG015zBpUHsGO6XFHo/KOF2t8jzTI2k8uD
Y4EgWhz8cFat3LrwO9QdcvFlgnkSh0U5I4wH4X9qnJe/bScQADidBiYWZI5Oh2CC
pgJbn2elCH06fcSp8HYRS6GPH/atMca1dGUnBT84O9iq/+aKVchI60ucSdqJdybr
MR+8DWS/6Ha7KBgVbVtC/DnCcKn7xjBC5L7HEvrEU15aaV9Ka2xqTGpQMRRIDSyy
mlhPdy0yBnROxTj4ZBHdNnZ9NEXnSxuMuLZbBuEtEHjo8pe0EOhHqPCHHrhYWh0Y
qL5XJOV56/RpSgdK/KJlLSl/rvlV0JdKB187lJu9sylLo/OgqWtxnyGR+zsfp896
JHR8jM/EcpCYqDX8O3HjKSdfYVJmKvFOe9ojKzYkVdWeC0pKbT87pacuucdFgr4O
siin0hTk9+qN0MAcAaH82NYkFjCnoArI9E3P3cOx1IqD7HZIhma1NMSgjs4PN7zI
9jITkaVBf/cQ0C66Tz/Qq8t1ABHFsgxNnPGrRiFgydaw63ZVpN93XcUCHayyEMBq
IkjGf0+sW0myzqnr6RJP9RK5eKVZvIBPkG2miQlgDgIKRv+kTZP/c3FLWaDfxy2J
qrPN79e62qqRhQ6QCGDM6nU6wFF7E7lMKhNPY2KKcNKG/TViMLdlufcnF1I2ieRI
yk8RYclaGsoI2DvJ4Uopl6dCmBV1qzhusukfBytUf0H7bixW9s9mSLd+PfE7+w1M
uH4c8RkkUY3GNNLt/rSc4Jbo9kg+eYJRbGSxBVuQ1Vras3LRC804u6Pg7l5G4fDU
UVZBc5i+GflWRyMAOX48fczLO893ndG4o0xzm/nl3dyu3yGUCyu5LGt3/PCFqFrM
8BTuA4cDkRWVvNgub0Z+/EA0ndM/0RAT3ZtFtSb9s34hbxWgxAn6xMf0EWrsOASd
7KscT7Yu46j5esM/DqfxqdU59L/xSrpf8aHtxMzyWaFJ5Z9y5Z5dI63o3K3VM/nZ
3JdMVg2aeLDssmGjgvwphQiq4TngqEsY8lU5oFkCNluX/37bSW3REnCkl1RDtFfr
h6PQvV4nnK69U6FbhR/QA9oHP8lOoDQ0dBOZC+I6kAv+irT1Im0OZjwFXer5OxLJ
EMJQuZMp4/SDmoLew+lKW4NwXozIE64rFWYbu1IhTckqkPi8IuFNP6kepnN0UTg5
67MF5raQQawSa7MayiDaNVa4tKA7eojS0ymKFvsysUtUznWzwyGbkkHXV0vWk6OZ
i2fGLnyfLgJKBpKmhrEjKOZigKbaCqcUhrDdwHXgS52Csu2XN53m7zkleX1wbOZr
8g9ZcnqXG27rghrUGN3Zy2HnHb/1+F0muLIAzxTrvRSQkuGVYtNfzBRGBYs8LCSG
4TTsuI8ZFQI/4/WSpYCWlqTBxquc8eSoSdcLOmvmWAG80+otouM2xG/zSmnKXtRe
76t+YoFACqoP3i2MWekkG7gT17SY2IwoQ2Q4UnQ5aPAqA3kzcSB/NWSAnSHenA61
KemCIJcz5tFfNYy8w4qRfNrMsDShIrs+0Sq+CK+N5/S5b5oRvw7mCI7GovGW5uUX
LXXrdkvEdIbPQdo7NptSprnjycePOSE1MXUS/LZTkKWTQai+DDP2keayaCK6nrzV
4CzN+FkjFkbQ5K3TAIjOV0AR2DKwQem1MAOJlYtcImQIAZAxDE2v+SaXkJhjgvwR
kqxf+gkOiSwLJ0t8vi+VrWioO+1pTJFvxsJMa1CNwYanEZCm1YFeDqmfQiXeX8/o
2NJu3fdU+Iw5BdDP4eNk7Mgkkrk4XU5H1zOg8Wp8zmaR/vsGm/hHy4RDzkv08BQh
0Ky/6TD8N99XlZVMGabMvPRQCDAKlnGH9145DSrpGFA1+zZlVF7fZWkkC3yxiuDw
CZXSQ8G9wD5oY6zK0VIryLWfSxNHTI9spoT2/7ByHBJDDtuI2W4Dm3E6Bfok9CfW
cJNwu/UjMNWzw7z01AXbl6EUcNWpTXPmVfVdIba/G47hyjRhXf3Yo03+E7m975JC
rNoHOt/LOJ6oxiuPKsB6ia2aedtpVzRpUne/5HQkZ+FDW98vx9bTc6P1vmpQUfVn
oNYRUsdCWlcenlPVAynkohkZeJZfjrxJ/NKQEyzUzILnFfAObeO6GdzxHLFHbs8J
ED3AWt76gtPPmnSxBYBtdAC9YYUnS2nV1+Di/1V0sser7oRCjsSk+amNUNrQjts+
ThG4YypyrOE3IigP8SeH6M1E1uc3eO1xoej6ERLWITbNYOwdnxxQK2AkdrzXi0wi
DKmdoVDYU+ZnFYonx3gjJv6IHRNafuMqQdwy1gLv8UeTQqeZasKb3XFciDY32cy+
Gkfr4wUZC63NsqBmDDT5AXHvIEiN/9z63yY109EO+HMDmlAN/2igoTkEef6YwYJl
LpZd3oBYPILdAHOs3Da662V4ZcjkL/2UxyP9CtPRKweFFdfqrTpmkk22inUDxKlg
jVmeX885NwGDuSszKsRpkbu2a6C03znEdEKOlk1dmtox46qdEnmmFbuGYVNE1JZY
z6oIcxNl/+nrDWCY86SZW8i9wRukZpTdvOmmLaz4OuOvmS6+wgz5gDzkMYN+eDDj
432WOmBAlsCSG3xro+4y4X237eSWXfOQnLWuUhgMKjR2b3H3kVjkgnczkrS7bpTB
vDE3FovqLgtKkMT9VDFv0CZj5PfdNTcomEq+9TE5aK+BtmmhIJfMdHjAGBM9Cq6Q
p4DdujVL/Qk2dYxkg2R0kLiF6sNRKzlHOTrXcwhaqgRSImuDiyZJslf6MvsXiDbL
MXTbdYPuzGsHmUaHMAno4G3CmvcLKPmoyoJo/KMP4gfhHHCDnqNdll2HWcr2Bv1S
tGdmwJDAE5ZkzxSxoibIp5HkdBnOBVyiJr+VP7qwSHK6N3Qd39n2z9gNGvQJVxVj
Mz9wXq1r1edCTOA6D+jtNFAtStGVnjIGsUcjMDLExa6L1tajGBeiZpi59mCoK+7c
MsuHtsxwAzW2DqAXwz/mekrzQz07CNyu7+Dr2nu3CjLUjRt1zfK5VtYFh0l6yg8B
lbV8VKDxw9VlfFbdetCqvpLdUCRziTzOCoPdyrUJxk+i4Q+agOoeTCGb0Z2izMAx
6hDlzmz+9RNCcQpOEGmARAcZl29+mCEyMNU+J9hDYzfC5j+d/6IDlngkRiFudx+N
M9N4GByfDOqsXpdqjHYz9sCdaOX0jLxPRwOjSUV4+Ud3mDerYimhkXU/zkM+/Jp7
phZ9p+08kECY+mq3U0ku/ZsErGe5O3slBrOIqVjP/C1BaP1GWFNR8FqFVvfOXIpL
Q+5ChQMi9uhJLagRruNm21VLrpHwl5Y9K1agyjkqNnc/LtjXmmhb6w9xhMVw1Ezn
zu/r1KvslqfLY0MRB8t0xkOCaqiHt2OxDS//+DRbhWdq3IJd8z4g/L7FNMtE+fmP
9H4f0wPpac5IeRSufDfg7VpCjCrUQdaCgSPbPeH92KepsEs4zRSf4hPeb0CPLHTl
DE+EcgyNIdPiNkI4qO7j6MYtku1QRLnuKPLxtnY9w1+IiEYBbMomR6imTCCowTya
GFYDhmH5276mbJPDUNkKo7m+59N3a15FNjL8jDTngzaSlUwnNwhqHFfgslkg93al
d2fJSjmgkh6pyCIPHHJLYhN3N/NTfBXADNujAHdgmkcn1xoCzotPj7saQjZSCVTY
QBM1lsfr5ilNBWTKOSx9Lo0mP8pVUkpE9yhwwCkmYdpuOfR41jKxRIU4eZKc8GkO
J2mmqE1PUbJzoIJcf6O/rwOQVzrehm9VZ6LnaRBcD2kdTOoKDiUKlXWWPS58bDCq
iagazYi90qmCATDJj4BfJZgRutM31wp61wHCRgylR84owJUp7/zRq/YO8dbSRBlM
oUcVuoG5jgMfShR1pLPAAVBioEMAIffsQ4akJPjBGf6/qBp2ThShchi6nGYY2IHW
GPML41U2yKeOYEg+KOp8mO6vkhrQEqxBqgJ6stZjXsf2UBXf21E1Smj1sQ5YKwT6
yUMWsWyqNw2fBCQgpeIe5A4rZpNlkJYrv89bPl/oqA1jI9KxcCC5+pqkOo1AtAZa
uXVaPqwuaNBqRibeA/5Iud2d22ydO0uwQgZoJgD57XL9zCyrxVkOZwSGWZfVDW9S
8V7MoNUC0bhK1lAPERpup3l5gYQQr6c4biLm1S+MZlv7YZdzUSHJ1w4yKQfayGKF
NXvl8vvuVwaamMZMV4UViSoNuRfJRSVKDJNmT+V7RPoJeP6lfZVYzJYRVRRwIW72
H4V35OqL3brZPD1N94xvKsNptlJolhGBXoL3+LxxM/I+BVVYc/30/VbagA8aQ95e
ObYBVmnrXmW19f8M6befBF/Pl0uH22N/WzjtjSDwZnYUeiu0sgD7Fvby1eoqPJNO
IXxrZGkTNTOB4r07fbOfj7gYSKiObbAEVrm/wxxku83cXD0oFlrKbdTKgj7Wz6Yy
oZDofzSFLeYZGouSmZ8+2HY9515ob1D+NU2gn5ZSE8v+fIpuQ8yajhHJ+L+fyVti
fSvYa5J4v59sIEQ4Q3IPMvUV9KoZBmq0gJHfiBTP/xXovART7UoELOL5R/0cXOqO
rqc6p7E/M0SIrI5KWpuQTsSQu859FHDkxLBRowA/x4E8Gbjft9RxsVs6si2XPrKT
D3f8XPVJemXVY9HUOkU0tN7B3i+VlphYf9EL3hrzE0EZ4jP28hh7+Kf4t5N9ieho
nNLodfN2zoRHaWQAnudUx5t+T4o9W4rICbl3k8tTe8LNAUIkJZxVnMA+iM1y2t28
h8sYVV3dpVvcC+z926yq16LX/qAzhWR/OGokUJWhWAkcMFOyvVmZEUx6YFRPYIOO
5U6XzXQC57VbZEIEpC6pU3OPo7KdV1s4UmEKmfI8xvOUMjMU4lUk0yGqZWKTvVF+
96BToMAlHri69zvwo5HeyKKkN97vtsb50DY/x775MviuzwBShaMb1qsPgGdRweH/
+t3e2hXPxB1mH5lCIdtC61apc73AIdCHDQy0WPukXWp3ARqYyfxNHHFFdJCQdPcF
rOmMP/vmm8cV3Swohi6FCa7as9fgLBadf80UVLkp3CEqM3OmOS2gTQ9+0z3MtVKT
mwRYL7h13Yz06DEOE2e8IjommkvuZoexcNwN4o8AYz+SO82Ls7NSWvZ2QpPmxGyW
mOA4YzB23/hcfGp4f0IJgkVEdWUkLuARpvI+wvy92prKYDxvu/rMLeJVB3I6Cf8K
aMVIQbdleOOPqw4W1eMur3toZQ5sRa1NoWAog1LQdO8hkJH0RDE+c0+ZazecTQhP
r3J/ZUaYq8ORgA+bRWXR5KTUqlg9HofmhtL5/MszO2pDX/6vao8e59jYtZA50aR8
POrBjS23Rjm+SHaK7AfK5QxT6p9fTWcBBPJ4ilF0HPhhFwvFnAuR9iLv1bAPMJlw
l5pTqsRTgQJ+9JdoQSSMTLRG+euVBsWXLoNND2l5YOIJo57EN0HRCiDq+DAVjfLM
QpNKOQ3t865En2MT6fA0//Mz15j0OQ92CmbwgPDCDSDgpJx3ch/6Cey23sRpAsZb
LTkA/iQVavtXMzSI2tUl0JuWVGkDywX8NbbxDeGFd/i86mNmUEYCAtQ1Z2UKVpQW
dQ/iC7fWFiMDxigEhR6ptgzGjhEB3Dgt+tfNPSUbuQ9vszyJ9kTsOY9M8DjGlAQr
KyYeCm6czlabHz3IRWGZ2pBS1q486tn3LpGVDAC4C6vXfc+ssjZmzrCfx/PNT6o5
5qOXsJRA1IBCv2q3u/toEFNHubEX3W0JUC4aUuDrr3yP70j3dnmIZTwoGF4ZPLAt
vFVgOH31ESWsco/iJD9GKA+Ne923WveckuTZRSJjVbUb3X9bxNTk1q5vO27Krkar
R69pyKdn7n8V8dmyF2I1lG92R2lBCNuYQIIHbA9+KETWyNvNi/3xWRKIlJgANhrH
f7qDbap49T+IkR8dBGZ9H+JcVgY6vtqZwggrlh2IJLoqUpjhDL9u8U8vNElsPke+
eOztR3WIVEG4ThjNscmo+/UydhmPb7pl47ecF3UU6vZmcBikIw9uuwWvyeeBkeWE
IeN3+hsx3dmGMVFP31DA8uV6l42nIeE19cSrkFTA7nJXdNHambtErlGZoRV6bif7
/XqU0j4FI0+K3Kdecs99XoadRBqTaNzeyUpxeUXS9st8MROoUQVfb+xxZ+xoxn/4
krtXJfpGc5o9ctihR1SxLx7z0Dh8uJPD9DRuhTpvFEFAkkpZ6c1fO9K7jqc9Xw4M
SpkimkZeIaq30vCkK0qU6nWcpKhFlFZKAxpyr88o7wxPmKofZQFH+MpCdalqM98z
tMCzGtvbxkrb3AcOTAhQTMwnHQWGkNjeEip8azz0W0YwErj1qn3KzTlDy2foTw/M
kQ3A0VeZxJTcvvv7MNcLlNDQ4CsdG/TCN6dYq9dFd9uk3M8QIPUwN1wgArKPbl0R
/hILR6MlsVaSVScpVyQH7dsa8x4d4j9rLr8WRKzYDpByjEuNocGua//d1EdqA5g/
pYthcHd4MgXrcj8BRKw2ZMMsyBGs2jFcJGAM4wyITcaEFlvR40k0HRrDwJjHREIO
GcW0fSgbrZolQqhVJjVlHdm72SKxcocmZ3Th0DLkVT9NpFHlAqg0QKl3C9TK2nI9
aZtMkvBeop2C4/fGVQUj9A78S7N70PPyqUMvCpyChUK6whE5NBwKVaAadZM+27GN
nBCUom5vCx7hevJp/Y20hDaSq+DKfTTMk9Ewy1472vRhkNDJkCi788iWWaEZDOPG
rd4juf8BOsc+bffg+HjRqwsZ0N3AbRNlyXrOnj0AOCMMuAd9TxlxnBtKjI3x/WX2
AnBDD4T1hLkK0Vb3fJQz5wntdz8oy0t+skNuQYWEYNLEJHX/d7oeaqSen/OiB2Gl
WMUQBpZJZeSuBfTWfSg+YCxp2aeSV10M/oy5h5IvRuDjsX16ulXDpwOP7cdmW5E7
N94qDcHJywAOf2ByKBO60Kq3ryCHLbVmaDu5/IJkGJD6vFhTrO0NukN/Ulh81KB5
KQM/2yBjtr6i+Jt19Vsumd6Zn9x7zTA4YsguloT2hp5i04SLa+fJccYOjAQ+YIoP
0GRtoNu+ja5i0SnH9wtPKCIm2/jp3pVvS7wE0bNjFSeRxW2b9VTFbmr6kIZ7+14t
uFEwwUNgcNPx7fk2mYGKiS5zTFvfUdAo+QnlEMguRI4q0A1eeCuYIzyNFJ4KoElW
8i3zkpZuzvtkmkAINpxbv5MNZ9ygYoDPGUKsBMHCl+NNoq5AY8w3BfHYeQxC+gAr
ipTdQjdpmtbtwJom1SFxFT+guMVT/S8C/f7aT52nY70XePEYBTyCfZF6ytsckTKa
pK4GvnchOtUjr6lCxos2JuwxQFuB3g+gOMg8pLCzICt86BEeBS0oJjCkgaZgrd/Y
YczoQdvrnA4443tW8gG16xo9eESbNmdKNW23JNW2DQRKy5anuPIWlweJD/mIcOrJ
3hhuUxSGm5N2eck57+G+LaapAsmXJm8iSaYgMYoolDE8EtXm7jRroCQASz9i92V1
Z1GgQv5T/WcSQ88X5l/Kub2I3vIfM4n21ioTM/b6M8l3YK8USqNdMGIhhJjQwVbd
NVPqcnyTIZlqomy1tK4rnj9BPMaQP3Ccaaq6MY9YpngbHAWnBhTlXpT05N46hCJt
is1b/ZS1fup5PirDpobYpSXhMOoo5tI1E4Gm8gx1418gtMNI7MWoZpOx18M+lonG
GHffcAZk3gidVqz+uUO8kL5Ze+VuT5mqhQZI4mvMvOnQxT6/6HrH0+z8Hnt9sblM
7Own88HBuPJhdffQNbXFhzsAyKANUv4GEPdjS2l28nUtuEXSubq6PUsl/Mk6GCQx
sphzD+jg1PB2uZ4/1kVXpAm2geeBFEU2WZ3+b3ryW3s2AfWma3vOUlmjbFTH15BQ
k3K08x6jvOcY7cullo3RxTYVkqVoqPFEvO0ug8CLXyC8eVOsVVYF9pY/+iDUFpNm
ixL+z4ydpsgL4IUYpcbsYj1Qm7S74zP1pu7lDaSU77yxJNJ44EtAg0uK67pN2KAQ
aiB5Xcm6bf3UDv/I3OcDcTx/SZHIxmocUzsQQuy5oQCjlrLJbMXo3a4rPVImnE+R
NqccTWMQ73HN8B/kMqrhdEQtENGt2Ra43pTbexUjGGgKb1+J2M1dCzjrE5mYY64o
mPUGnDJRHO2Vw6Xyw0xQ4coN2Ikc6qiacqEd5w9dD8QoWsrH0oyMlIfPkwYv7/EY
/4XvGjwuILkBJMXm4ZKN6NKkK5KY2LgmcK7oKedFXuiKFJ5DFB3yP2PMJv85k9l8
BbUfKOJlfE80/eRxvx2xYrRAE102mfPcZpDOEjnSSdO6YjqcYgXdAhuOE1B4j2O2
s7ZuI+4hP7B8ikmQ3QsqTs90DaJUU/4Pdr7r7oRg4RBYIzUtTlEqlUxSeqi0qmvC
oh4oj7nykzdEYM45hyVcDzbD/6gu5Td1HxW06pgQv3lG3Kre4/QjCmUsGx9tCyY/
EKS+NxkMJh4pUciXkwdFs1htcaQQ6b35zXh07tznbejv+BDBfr77+F4kBuSvelTD
GPAlB0kTA22fsQpeB5rXaZT3cT9uUDzP7Ez79caR4xIbsVixDQDBDR85D+4IwQmD
GcPmpCOXbwY+RO5I0ZvEDQhA1Nm64iCwJ1UKdvEhjZ82zgJmxjBS+OBKkzjqtqGC
4e7QGG3rEvX1OsGcCdF4UtPGB80P2wszKtxeIEcGjqwxKiR7RJz1DqopZ9V1LcdS
jRDUHMZTCnOHgYOtVUQuvxLo9BPvr/q/7rJa3z8wlxja69ogEQ8/FZosKIBALyxU
J6/Lxh09AKbfGtUbwhG9JNR+VmDIw8Tm89ZBE9AjVVdcPlRu07Ec1hxEOUnxr6oq
ARJGVT33jHmJSRd76KDHSCGWWTEG4ev2PPmvTYlElfInqOVf94WSlEID37K5dJwn
Eby42DjB+7BE9ql3OXDfZ5jFRBZsM1bA1ve0Z8Zo7ScefUEn4QI6pMho46G7lHQ7
4r39p+NCJ8vZ+vWj54dAPZcg3BYZJKoCsZWg5DAjzd/e1NTYhPpa0aHuTVOHXWBK
xnUsrd7dD/d2d+/zXyrkEzvxbFed4nTtTq4WKNDyRsYfKgSIRK3jKFaPy9vjiCNR
1ivzXEEbNM+GZYG79OfW5UGVPYWBmfKnO8sP9J/wykYvmSIrgw5jCWX0qT61yR2e
GBqNgg1+sRy/iROTrF/GUGWcKQwxmWM1AoBsdbmIkyPtWeMFY4HmCFyY8mWPQ4+6
LT2MZxr+1YszJo4QcGZfVGgG6QkAs70MdlvClF8ANi6/tHKemfiKlpmQNo12Oj3K
VD4e3Z2q1RhyYhUSIxZfZPweMY8R4r/teMTmrLaRkgwJQJmR+kYxkLPu+CP8f/m3
YDckEo6qzr0/n3PziSvdoSOxC8OxQVaJkrX7qHzerE4XGPR90SQo2PluT5zRGyf2
2Hy9hXfdlUtxRsTcNrC3g2ZaemVzgbGmN/JLrMskANTLWkLpEzwNH4UFoJnc0oZa
YSQO26fGuQI81GMaf+VM6WgY9NHerWwRtkS+8w5GMAWAu5Dt62RUJDlfUEreOr+U
oBzQWG5GfKdjnDo5XmTkbw73VthSsALXmFBdfpclG86mc/cI5XVrsM3J3ULeIpqv
jx88wBYpsQQkpFgkN1n54tJRRyqM3cWnbaqahj9fKOMxfNxq3dPTr2nAbIJfwzxM
3M02NQ6gb8GUZR6cnERA0yZb9MH1tntXmvAf2hWfW6wdJ47Pt/heg93H1f7BLrMk
2XFxkYaWfOEOWO263fwuwc933D2/ZpO/iLTFYwb2/n9iy4q956iflRzmjuWYyukb
IQafgnzTt03/Nnmfn/gK++0E77WZhLPTG7qj0bnjrnH41RYMNl2FiKJGRvMrkkJ2
Bs8YoVx/yj8tDul1eSqNsUgx0xmMCk4r+/yB5nzB3XvZREoYn09W98RYi1wflgBd
CDg9VxABIYoYVnoH5yt9/jmI36RkvTJbF69uXt5wkyuOZu6G4+9Gu+opT+NuFx/o
zj/4yoVAhCUadcOqr572sRZE7fqInJUXcfXXt/T91uwZFE2hpQTsKysBGRoQ5weh
m3e7OKwUuYVYxNjGqo5XBytaLTFAFRYEo6q4lX/K+aSbP6UoZzC+mEGGOVLLX9Tc
5+z+rla3gUZ6FI6VBXHMQZGg65AfQG5aNcyK2BXqcQ+8m+cmr3HwaBETARTMZ7Ap
LVgcEiB9Hvb70fwpF0Y3Pt653VyU7CMuPEtqwOsoDPdQy1rrI4vMS8kyVY8pM6t7
5GW7icHrcJeXuPTUzICNW8sgbZYLfDu+75gj/ai8+PrUigUWuNCbN3KO4vS3X5WK
kue4IC7DvRUVUQrF5J4Hlx4vnhTv1oNukaPNcKd1KPfBxfdWC3f1uQ9BWowHY2HG
XuUueih5jlxLvwe4MksEdDK9pKEHV1TLhzIjaqhllFyy7WXiVr2/xxPYGUHPON6E
xTDMUxYqyHfb0AZwXqTFpjUQ28qSMzkdVH7qJUeZrtgBiknTHruyB0//ceB3PTXW
TScLtcUg9X4gU7pU6glx+B4kPua8r6G8nuULx4fLqlnkK+iseQ7JJ1+WLiEfSxRc
wl6Ik3yTn1eAcN0nRWPRAXrwYIxLmN6SGCQRJr/SG/lt2NG6KZs/y0zYGO1s0gK/
vvc6XTbYwctzOeSbI8EeRJcE3ZKzNKoxPDo+3WTYsRGPCrNepsgFWTv8CkfNUUee
0NWKl1nyPheSebXUGpomuNzKSXQMf6cqIRrfj9knUagB9RrPslMvPCQEI8Up9xZK
+rQLdlOI6Bm3Mkhmn+rhsh0XsInx6SXGWnOLIfL2AmITkaHe9VCaqbjNsr7iP+KG
FmDBkgy8kBqPjK1tHWrllf93MxTPSYq8c4CYQEH50v7hBvrHm9vdgUV3ouSew7m7
YipoS7Wh/0jb95Ojg2zAcmR0eXZRgSgUXidisIV9mmahaTGGV6enPg5RoEie1sw1
YZOQhCXwa6VpyVDOAJnAU7JNd/fSFFr5SekStZ0esmBH4qa8WremJ6wpAqGvMBGW
yKmj/cWqP5y/LIZp5W8zd9UOm6AkOHyw3BK/xa3OhvUsuBURaS0Jl4W3QdqkATwu
YPueeEA+Gx93MwTHMOqvmg4DaWkMg0RaqNI5RFXG+GyvDeR0ALVwFnmfaFaYLADu
fEoZag7nVs/OzYcpcQ3enOe6SIyk0ClLA+kzp+Uo3doUv7qQB2ducxMbnhkUTJqW
FzVNpJQQ9TG/J3lPJADmQYvyjMLnDx+GwLrDM0W15n6Z4hVHz8M+FjCqeDYJu2tb
ySjFv8DtvbsV2PvqBfTORLg57xO7wTc5QxUAulEMObUw2LT6m0L4ulwwH+WLgfuM
nLBcjYUCO093UBhAiBAISkEYPlmxQA3MuBcgFedvxKehKL95Y2alF3gqFWXGj1iz
WIenq/X0BH0vvl/GsKQBPxncp6doNvD3ZtIjKGqm7mgiCcvK81totwzxFYzjfYv8
1yhQxchsAfiS2IWR0Jt0/5obK1lC7mp/gG4aIGFLCSTabTfoAgtkR4mvwgFfd4uQ
1b+v75HKmmliBsfOydtmFhvOjSlfVuymmJpCKZveyVsNtU6P22flzfiDz0P1bXGa
jUHgt/zmOH4gLqdE47MZnU3IbvXXh1nJ6G0+CFY17RJezm+1hwALtmo+D41/eoK7
PcBNBWmdMevBwTFr4lHgv77WixFJof8PTrxxPxWlZCYuUsbojFRUyD9soNoAmQRf
nCXsxwqW8a1YQ071fPEmX/nC8lRYPG6V9cStMZFPgzfOz6F4jBMheVudpYRc+lOK
ZHB+5UcDDB2bOTB048JNfJRCPPCBVs+v7m2jmOTQRkF5+vG+dZHrcZxQmCgLfwGf
4GQPbyNXTScYrMwahrVZKsSMX8q+MeVrpDEfelYXbF/Amz2A5q64gNY67eRPYoCc
Acjptv6JMB3hurBpo3bgDyBIx1vdD4H3/7gydCBgfeMXtc/JY78+qTGJjYBXI6b0
o+LQdGazfVz/++1ZOjRpP8+XfJFHWw7FQ4bGE//tMiDuyXemc9FfkP8OGsety8X8
gPRXDEuLR3pQpCge1c8Sx5jcPzm4lnnDwnkhwpBApP8fZJIw35IhPS236Z1v3FuK
E9inB2ewRQelWKvAfdC11qR6uRQmq0xLKwMlVqxQJ5sAEnS7lWghVD2kuS4hfh67
U4EXm/Az0zSu490n8Eg3Ql4jLXutvP677UQgkFVwIF8ZWArGxLtiWhLtphO3X5bS
kMJQ6ikK9U+IcS2uK7ligUU0ymt8sj6GAJNtG5A7u8532Ck7msMxZ29Ho6CATl79
HZisfdy1FmxgDhUQ7s0+bcxaKqGZaOoI54jrT+A8ruGRWQAlbFMA2YNX/RPR14YV
7pGrFV+imcxE1S+ezCLQ75HyJs7GDYQrKUIP2FoTUYkJyXTXcSSmzU+T7Gkqzlpx
EaYqm9s3sIaFaCm3MVutXx6JbQxN+qpk67/j7CzI3hZ6ZE3D4+Js10s6b+ONC0p/
5EkZ9Zw8d4o1Tp4h95e4YIRXYGZx/rDTtYijHzmQoj1pPKkMkyM2F1fZtgZsjqIF
9Bv2lUsEMhAZKVoubgvdXYqsGPE7eCfOsAj19KhPhd24pKXPMLhn+9TlPOKU836j
IOogTU7YukA/9egcjaCo9bRs9UKECf01JRJPlgnc4TIXfZ3lKHoQjk/4jre+8Hul
khsBdd2gmQNiZ/C3XCPEMm8LpsEaFMzgxcEdg9/qL75+5S12ewEtxQK4R3/RKkP/
dRbHB6bE/80MYmPMXhF2X4eskvy5NDcrkZRTMO3cbgS472JcLK+wnTGDrAIFQjbp
Wz8bVD2hTTstcWjWVKLssAH2RnTAch7zSVQWHv5awmHONRC9s0RnBYbfsFtifeAd
5h2SQ1bDlJQJr2QKpUWk2CcHwNgj73j9WKYbpUte3CFbofK17w6r48s9O1igomm6
r2Luw40KYFDgPWpLTcZlqBV5bdkfIIsqbAM1AO2FtDYm09Px+HLjObSowdRDpOst
L55lvU+Zu4OAvUPNGLu4PpRLjSORJKelIzRZaJFEDNM1qpSdOT3d82GT6SIxPKEO
h8B0PAp1LZyP8oDkXXkCiniw3AmReieGqrJ3F04xXkOZO/wMK7Rag1snJ74Ebhg2
9mMHDa2WQB/58yb3Jc8etU1mz+4s80TBFsQ3sDJhtjtMLUtD0cTduhJQ+c44AHPx
VVID+J/ka9BijVQAEvaO6F71ypfHkp6m7hhwz1n9qyvmA6oXf6c7PWOEMy7Y228T
kkpyOK3qz4HlJUZ+n7oP+mr+QJNPR6bwyXzddBrc5sVsoeYxCk5nDJxHn/UdXoAa
CmF0KLty/ash/ez10HIVIvFWzKObFHdkkdXqUHdObKE57SizhALpjKY/8qC101Bq
j2HopC/kMyI/AS73ia5IaH2dvEwWgZSjEv1zzwFcTjqgB4AHzD90xDU5i/m8YLrO
aDd3KBdO+K6RTS4IkbzLi1jkR9WOBcL7cb/b9GObk2UKXl0BhGR2bNrkiXaNCoYN
D585UcxvYkatOEknaGLkwAaZTF+eglsmjQ6s82yLXNT45d/QWMMFJmNON8AxyXnL
U7qCe7yl33CGO5NlRISUvM4SP1Yc/gP8qRhR0PXV2Dw0YP2bitZGMaAqb/P6g4lo
KmTCrKr4+O5Oq62C0+W4xWRlxnCkup1n1cj6u1nTJ+1Y4HCbhQMXVVIecWg7d85B
poN6SC8HgFZjSrlsEA6RZgckqP43Bz9IHvkAkKDVxGJ2cyTIZhQKBRE288oy4XPj
/eGrkn7ZX1KxF9Fgnqqkn22eH5d3i2NetwauNL8RZArqUgfK96tFkWD8KYgS3bkK
8e7oTSVImDehxECS4BwlY/XZgks9QK6IXQnADaozPaa9UZgqPGMyaKLKZPmSgjb2
2yoJXDnez1lH+TVUGLFDio10g8exzoax10st+R0kK+EmWT49snsr2Zv4GiR+Lx0E
jxy1ocaec+flBhaHxWALtYsOvs/Lc/BFoidcupWqrR4yr5akqjfkbQTkh/gOliP1
gUXHlgPD88PYwpWL9kQTZzyfB2TiOsyQNKfheQas03ohYToL7jWQhyitjb+O4Qtv
jiiR8jiS1wIw5AuWiE6NSYj7rLvA77cT+X+uflDZraq3qpI6RD2lB/KuFAY00cr5
VaDmEHOzEhhy1/MifsZXiKHnq48R4NDH56wJ46uV+3Mf2RZ2WyStPdSs6OjXcZM6
NOd7v5CfLb3FypmSTXJVeait6nmpgPIaS++tE8RKuSRm0gfFSZ3HMjfB5k7wIy2K
HnlPsxZSjz06G6PGlVXeEwlRttSftdBZCK6jksoQOpkT+SQxcL6XBBEuh6P8FZ1l
smjBU7kRq6VmSA41e3kA7rea397zil7gUEOAQrGUMReF4Uu+N1o1DWRAJk8bHFA6
8/e4ry3fjqj0RcqLSeOnofWE/jX3WcX3E+Bhz+2OkwtYlK+AHc6wdBzx3F6BEOTO
rXGqG8HL9h0MgJXBRBDmRmdfjKjE+J7mgnUSXzhwe5uxSb8FtTLRvrm9uGEzzmq5
ZauDHABI1riDKudm8F2YwTdgJF6KAs6P+v2G3BoAF5TXPTdFYSbZIkXEnW+OBWq2
GhmAyDWhB3xCI0cd4nRvotrqVIkE5in0ENAhdJwBjSQkPoVuyWvoeOCvYU3iIWo/
h1LUzjxvgn16jne1KRYDGU/t6wt3sl90Kl9yl8T9xVjZCXrzUqoYtgMyit4iPipl
5ESHVMuI0n7lCsy5hGRxHxgZg36QYADDLiGv+FFY1lYFjxzaXu8p0oHpRMx4T8ws
QLcCotSilyW718gjcHQuwNt+IHyD4ZZ3k57XSjXqtfEqwY/4+kJHe0oeEnw3AEd/
csXYuVFIbq5wcg+XsTMrqk8Dan1tVJT7njpabiPo7WpuiUW+MW3SbuOGW6SxpN/I
7aQO9UDTxBtQwrDX2KS1F/ZfpmcOQGeKWd/Utlnsb9rg/PIv/bEbYebhSFHKhh1I
Ag1sntIgDfsbZLwImDHpgm9wjs/Oq4GocNkO7tc1uxqCS67M9XconyzW/DTxgU8p
+kc1B9gwBw70w+8SPRVncZ7dgmZ41OThRV/y1sdWfILlaOJ+3OjXGJqWSDnfOd5D
tJ0dlUe57pWDtmCDOwoH5DnbAOZLSvt0QTXDhUPmXxU+SbyxEftotvx3+6l1ipRH
7CfXLton4jbFaOta9e5ZkfjbigCqrAqJse0yhvEn7xBvdg59gbWpsy5j/I9O1sNP
ncdcyXndwiW3p0eMKXZAvutjErH7VDILgAfVO3JoulLIrAce8x5+Rc4HENPO8J61
K15zJ5IJEVmYuWHWB4D/d/uv4fDublMI45Jio5FhNpzgbQZl0O36L8Zb+9BXtd3v
7I7wTwaY3AJxA9Wz6Yyc4OPX6eL8m8AkqtvQI7uwDMjnajGxC3APSrZwXB2N96eP
O3qDCa+3kZuE72hBGmLdlRjrjfHZwdjxw7Oxk7X0Ylg8YZxKoc6WincmfqE17ogt
LU4xw20YCGn8ey83OFZnhVPJHPqxTtLY4yO9DQhBSl+F21n1dJjcs0jLfaj08+80
an2d/xjvQKhoZfKyOtSkCm5Hf2ub+dgijYamEjqNSIknUMwnnRAkODiTDiSssR5d
uxOx7lNdSXl45X19Z8czmQdzqD0V+eC+X+yGv9LWPu9uaapuJ5TCK48eI7ZNerkb
s8YeOGh7IEKkMJtVgVkZxtUl5WEYcXqaxMKDhIKHSOKWW9VEzRpe/DF3Mm8xGdSr
2v4yEvXXzNIA6hI+HQ66tO/ANaBd3I2SKYYaSAyDU0wcEnkeHxvfQF1XrbiAYPEw
fnrrMLHif/2aCpVFH9OXMh6TUDVk10y8E/qNiuCXG+ct99p2uyLHUAmiTQA5Ipuw
9zblCIn3KSkT12AnYNlTcWErRcJ8fkRdAmIoZVumoaB8nY8Di0kMlX1RKJlyUJ3a
5TV7ppObRUNvKLQv1j9OZn4WZiLpl6sLuZ9v6ewH/K8cIXBC2TAKznRYbK8DWOHQ
DbaJqy/grqhM9ciR2CZXOSPkXLAVgicCcjEElm4IQVbz6Kk8BTZoUfiK+z9v0K04
zxN2OBd55IhYTYMrpFoGNx8inAbih9UqKXx1p3tRr58wVB7HVq6lu0+zlE5TvV/e
AvP0Q/ncgJlXxmJ0OK9+0NRG6KCkL5OP1Q0/uXz8xciK4U9NMxgpfaqem6VUkNzn
h7Tk/42YM7if0LgYkY06isUtd707xgWaSWA2fcfHc0YvRYa80BW4FSPzdlApS7Wo
rmFx+BkNnC760YE72s7nz8mNyTqM1uztMFlPt32s+ukp67vcCrVdqyvo7thz+i0Q
rlreMlhU5T2tzqOrbf343lLvRMwn7ouv2E1n0UtUfyVRGgB2FIytvHTpCgLY9JV0
tPLkV7meh7EtzuUlO8txyI6Fwxj5qGOqjqYUi6zo02whnpqlA9vK5NDhI8Q6b/nh
EuwPmuC9UBRGTQFAEKqWzEFMo4he+8yc2XoLfC9tz7+nUsKorDtFdueFFBQq5OgR
Q4GbjwQk5fRC/d9fiYt/s9vT+8tMt4EeD4fL12w08ni0DDfVftE7SB4MC5ESggee
CAg65COqrfIM0BW+SkolGjaFrrl855uzaH8Ro6Rf3F34ja0rZGC5kImgOjCrnZSW
W2IAjfIuxzSAnlfcdHgqVOn8M+iGXyL2hH2Qd0MHGzQFTtQgpVETiW2RFGmpWB9W
yi/phmBjdatDs7sPf1YM9TkautbeBgAMryU7f0UkNSuHrTcoTotMVyZfQr1lb24G
aCxxQWfnKLGTPP2jJrkvWIW9Ed1Ml6gR1iWm0/CW08YJrSTMKuSOLrlotKb0ZAow
5iW8pIS8Cf3mg62Wkw4X19UWbvF4zBYCmdabXU+yyaanGQovXd0+YmhwcTsfrseT
0mWY888U7A1PdBuvyWPoO2B+d4kUbdI1E2Rp8BxC9XlDGhWpc2h5/Ax3vVa2lplf
1lQcAKrLniLSVO5tHR0EUEjvgxpKIjpWLQBQMlt4Riv9YqlnodsbZwQCRaBBCK2z
4dVCSZ2Jvqp3erSBuI/pO/bpKtLtjZrOQ7VOFtoTpo3WMBSEc/v3tZmU6cHidhIR
jqu8YcnBa7knjgSBAwrwAHdSV2FHEtyyJIZ7CHQGqLJ70z3rAU6bunfcMVgLNqZ5
/4VAoC6FXHto7GXoGxeSx+4YOLNNS1d0FL7UdFfp1zSJ95LFeS7KMiYQttcr16Qq
oB0+u55nWGR0kJlJzsfAFAKz63ZGEqXNA91FDdIAhpTcfKeJgBusFp5kkAmowkwb
dVMvEyAftyn5ZjQsVEmKXvsv+G+pTsK0qkf6PWOa0PjZxlzISbqTJ4e5mM1Ur0We
RFy2dwIWgA4NlNsKDCaLq4XrvTLJEuFm3raZyGhacPLXxuBtQgrIiZ1TjJgOqf+2
efwrJ6vaSIDleI4xqaBikleICK+KfnpBXB+zCAK/p6RwQ37p6kjgBWhx92IRZTHE
yayaBENEFKlvjv0tYXgMr8C7aXw37z+E3VZbF3jL/KqAlS7nKruBKVrH/qDdHpuR
sRQsa+WupV9aXnLPnLwFBls4cyAF08Gd8UwMYyu+LJXZ727zDsjx0UCW/5/J80X5
dEKc/XNyk86A5Pe07b8xA+KJwplsI1OJpQs9fZEBItI0mZnoc9+aPhIVbhp38wxb
7xBi2D9TwlB657TCx35gGni9y9GnBDuEEHxqkc69cYAtQgZ2ooG9zsPOM1PZaymF
Ra/3UeT4a1QQd2P57WiLYSx6Yvd/ZwoiZZYnVeA//i0OcVtQpJxsxd4Kji8Fmmui
LPmjadSSpSBfzebV+EAwMGmgBoyr4xC4kdrrSGDDItHJEIUZZs9evaIjaz3RK8r3
+WDXYQt6/CfBJSXq+YwS3x1RctdVPD+fY5/xp1LRD+LY6POrjCLSCiuCNTHktiJt
GAIpvy8LteYW/BRq/NDVeZrJrcXvOD2WxrL5gCDX7GZDTz/pdWApXO48EkK3kqsQ
raf4l+BLhNfAuJLR0qTZHurLLPMoIu49pN/m4bE9nQXBXm/3WVtYKvJrZ5E9I/v6
E9yBylDI+nw7DAMqz1iWAq0RgwgoptPd352MfeCduV6/BOCnW8OQwl7EKDrmPVjL
w2Obz7Hmf1lO8c2enclxHMwvmFI9ZUhewPPTjwLYxnxic95AIpJkMsxiPQ7n48dz
4jAX8mG19SBhSx5h1roqO7ouBL9CV0nXxfkB+QuMX9PzVg+EKc4J84wKQUbqdJdT
6EbHxdPg87xU3fN0Hgij+2jDB3b/u6wbYaJPk5eMJGCGY7V9k13iuA68bON2tij+
tX6GlxpsIMhChSvl0SbFPp+TC1lEZS1aOUOGiMn1YW8DRGMIl8dPP3uFklnuPDwK
KnAB9UaIcSRT1uei8Qlh7SvXMgYfUebSEM4egb6FGLmtxoFDqbiN0KApUuHvVq+Q
UAcPq7ZbkdTcSzEumI+guYM35HaHlG7ZSqVXgIlmYRyzSE7zh35jgyz7386/Tb+7
zc2uEeKNYXb3uLdacDDXQEUY/GTWIxtUadC4iGT4wFLaUiCocNjyJq0RS4evcddc
xx+Camctv6TqgEaY7MnEHE1c63t1yvUVod12gwcm/L5xGCxZc0GY9Hx3S9XdRuFi
cs5otFpPb4YFLv31/aR60H7HuYO1gydOZYeqGvA/t0VEdDwOqkYkHZXfggCpy/D7
ZjpQ1EvQbg8FVeL3hYcAlKQlqmJibQn4XwLaAsQDjprlx/XRnKaWOYHvuk6H9rWP
5ezgPFhpW7FCFXs0L7+5tr7aWrcKFIAGXItM0RWhZHCc8mXF3KtFQq+XYVC5sLw4
d/mO84blRcvpzMs1pfE7PkBoHD7ogP51dzqLkse4vfUQpLAodwoWapCfxfLQ9H7k
VpF3k+9qnoY6nDlDg2XBY7bJzSdDYLI6eENECn3/wmMBpP1Csvps0HxqpBkYewIN
dGMNPqsGSjpLnRGRQmq1ga82/kY5brucF2ZX6QLk+d+8EOzivKVI38rdwXL8i9c+
pxrZ0X9/Kr2jYSVD7z+fZsZq7sEk57XoDeg/6lj1S1Yy23XznB3Rn+M1ROyrRdmB
WxLnzDJiVerJOiDEGJsUvueY9oBHGmOR4IrBX4I+cAxeLFpKVCFcHvym9qQ6NRVc
+YtCjdT/XAYKqWleRXg48+fjedfey832xTHahfq8OlLZ4rEFBjjLGFsqjKwas/rC
vXigJV4jBzyL1FOu8sCTnBjgzfH0uqupb2wk1Om0+IoaUdGJaNGUYKV2bKTmnFGl
5dh1YOpHtiez9xnMWxXnKiQ99pSLc4oava3vinlT8mNn3IM3Nm+3/NW5sNyZYvjg
tWsZaPPUUf4Ps1sFd1BTzXpX0lEgc3rElcwty4IsdhWFF/JiTD7aVob/L/H89gQM
CuW/YbW9iFIn2aPIJolMEDzk4E8NFzVruHDdFQQeTYC2WjrdABYlqQqwJ4IcEbqw
Ma0iXkrOVsI8l2hWBQQDGAojN7qoO3IukkSHjbsiJlLVvxScOGMv1VmqeCp9slgF
tjf/+QiKknyg6O0HHSApoh/7htvG0hb/hqtC/rfXqxpy+b1oy2uUtL21OE2oRKw+
ZP2LUM133cal5ovY6mocPUyTvluHCshQMoRPlw7TcyAB98KsuLm/xFVnelcIPPLD
XG0ckDu3fdfPBs9piH1ZBBmly6jg7w0dlQbG0VKrfzft8J6toVm8uk/CABBaD1vN
vIEMBhxLEDPNmtAkF1j443N2GmbMd8OFPgPqhfb+z65CWqlr1PvS62WynOEWcvhW
Ww2vCgplpaCZXcOSKR4Tvqy38SnXuckAPgf47l9qAQbGNG631zqlhpNGvtBy0mFK
clrkcDj+hkbyQblOZAfF3sRxlJed6/pJ/zalZkSppfD9UG+9BND9tUZHCdy7i7yd
FX6nCwe8N4faI2SwHuSsHODcv1sp3V9V7P1w+aljSMGv+LdHhqmhveJ9CxQwW8DY
fmB7CFfCgfT+GQhemOfPdMGCDh4LulEB9QAKl3okFjJEaouDj2rMQYGazjXvtTbD
CaZ1/0n7T3QmoIR7uK6qPvBBtycYtDTToFMqyfk2SHFS2oGptk0Q9QjRvdDRvX7n
H3FefxjVWz8vGPyhEhNBfKWfiM+jV0UaHSK4opWvqPdAJTOu1j9fl2QuY21dkKIH
O+s71lnN+nydf1YISlyi4wlzNg31WrmT1cmtfPAhCjIefkr76OlKiQ+Wf/CN45lv
amV7o9xJO3zWBG0otR7a9P4LI/UIp6jeoVXYf6hHgzbfnnuQ4IYLTaeGuTIS25fO
QyWlBccl6ZbnHy/X263VN5JbHgwhpAVo+WcVQPcFrKx0sXTl+jabFMxQkR3kQXcq
b3HvAzlGAw3fZBy7u/JSTANHUez12npvQY7kDAl5xNJuQqNUXFaRElv1wjkyqly6
hDcovp9+piVEe8MuU3kNFwkQ5VuB4yCz/S3QBhQ1xMiKiO64pFcp3W7dXRmNabkC
gfkqm5Yl3T4OjbKFBGBzYpPDQEIvZCLwD09mywaE3Fq7Sysk9kRgcUToHauWWYeN
534Hnz3NmjMDE9NXUzWCChBGlu9F1MwIvKqauZDIVMt39xmjsqOKa+3Kk2MlAMza
wN9cuK1fO5hY88pFjh978+1an8j8arUgDrL+B+N4jrtrfgoBtIHCXkU7XK+/rz+M
mY7FYJpp3ksH8lhF6KgkAN5Ubu0XWEp4YnTFgYedq7nC97w89WRc1ayFqIFUgIkz
QF562h6cWaiGm3UZvsi8NUcGVcLAVA6jQZZjt4FGEPNLzuAmx+TUJ5ZkqgFGkH30
H8KN7XTPe+ZcuZEzV2wVk8IQ7qELZCw2uQ8VCclVtSzbXD6jZfIaKvjYrkwYjtMa
KrOHFDAR4a2rDHfp7NeTuxVyxF/BTrVL07Qj0+XD37vFKbgUeeLLtBX7RUjNZHx0
CKA+hbDfYEhEBjhjOeVYmH1cynjuLIiAd0UfJh+PNE7o/mowdQvBMqkRHWq4asRE
EhHM/1PsH9vw4Ud99/9zRxGBcmL+7KGusUgTHERT+xqRSRpyC4FvYljZr0QSAijo
cGDiup9heVeDKI8TmNkYVlfxgXpce+6VVU2ShEqQUyOF6dGlh/oU+sN1T2/0MbBf
7M4iXmirHoXWfxm6r9A/u2Yvz9XfZRotIRIEBag9CIWonqQZEl6kbXJvEHrpG/TF
6ZWkQsVGFf1dyG3DppNoI/YW/3KF4bbBEdIt1HbZfeGECUb5XWPDFxiXU6RGFGPf
w3l7LVU/SF6uYCxVuf2vTWSUpNm+MqFwRiANesKKdzOrrKU7Rt96kuOjxenczosO
TKzZ7GRyQh6fhCCojdeLKWQEEND0kMHHUIEnfIst4RNuJBvM9jCBHJfGzocplDAG
Vdl75xmnWRhfltdiIdtNVjSmoXpHh1hpafrhvN9uYJDhS/xu6Nb3HxkCwdGVBLbL
PPSvOI+IE87ltOtfBGlrfI0lAsP8EZue24Me9iQmEsW7QnGT6UYBK4aKpAy+oQ1X
Ewc7eGmpojpqey9hFqmKpPNXCwOJ4dmL3INnUFol55iudERKFBm+9vY6CTdvVigO
kKcLkuALccywyG/aZCudRmlfk/tcg5vhlergVx6Goo4SWR/97zwxi1O/dVKOtPH2
IkEgMcr8qD4eUbqvydyaD1u6lIZNVHTLaSnyMlpvTpf8U/L/ooyWif0ye8ZTOAmF
/CGdomQWMi0pArk4kL95CQciauaeceX4ULkbqK/Qi9VP3zrdjdaSg4ue8UhqDzmH
7hBu4ge5LsQrMoR5MDMZGKx3VL5adUORBzTHZtNFxNCvwD6BFH56TkHt5fWzerQK
WV7WW6vgn9cc3+tee8YhrXOmSBY6hCkpoMJCpFvagZW9ee5XQkOwt9IaxH3sDH4w
HassIswBYsPkvFNV/sZlXsBc3nUcr6uZhiE4sXsg8zqa9KE8+2MTZ/VAmdGqBRRd
rjiUGS89B1CWtYFX2N1ajTXkie/Ume1Z7hStTS11wUeLyhk2ucr2SNiHgwf64ecL
Lk81gFYwIEYUOs7jJfJi547F8kinhB5bnzad7AG59qtay5YbXlyxnkdCAyP6S+hG
1ui22Sly/6enuGrZSxQ5cfWyOZookdeQ/t1K481hfneE5fWa4jD55kHo/j2gJXc9
gKU5s7GUGMOlGl8cYIkNCPwisRRt4tUyGseictieBl6cZnYhTOxEITumJL2oaiIY
ZIDsuae+IEmSo/0nH4VErkKX+L7vRPKonJ/okGCYeL/mGRy0H5mXwbw0uu7yHoq+
uz6FXYznarA8yuuBlMRjO7Wj3Orx3wy83AhTyB5sIIfAxlVzsziYRlczMeps3X01
da1IvmrviFSi+I0WjWEY3Z/R6eXjwtiJnUG8CE2jtyfU0Knpumyyyn+5awBNKNcs
C7wdzYeFRF5PnDYGGqg2awV4+MZ2qJOfBEQCO8jjDdqMlfpc5ryw8MGGCHqfilF0
diNV9TQ0NRLJ53SynGXCo52lhOCDMjhdm9jrC1nUVGnGpi2OuwaHCeCCBjUr6eMP
2SwluybxR0Hf9T6c3Qg+wp+aXz/G54O8Va9mdyJmF7CsO/pMOvDgharVi5yXczjI
rpl63L9vpsAkdZ9l9nbjyFrJWIe5ZdRfT0mgC9TODC7268BcMKMaUbUDzVHtnIAF
wnMZsefZNfoOEO5aSIxd30Nxr4GOF6ssn71bUTsWOScon9ix161lWaKqdQB0v6l7
1fcdxOUdzKu8ezrpaH63GKS5ffXUFB3JtevRK2O5Ww+nMpJWIf+vgGTEUJfgorF1
3sCBTHRG66LENBbhFM4u+v8Uy5QxZs2aCgdJXgTlVNv+Kbo2pK6JpwRB3gBdGtG4
FFrSKaDg6Q4cXroerUfo4hc1+REGYHDlaaaYB8xh+hAmKrV++iTl+RvDB6Cj1yHN
Y4BWVRcOFAdsdr/8sFCcNQ3Ib5PMb+dChjXuVedkqJI8YclWk5J8x7kMbaE07av3
IrI+9GBE7hDXJJ3pfGd6CsvxsVYcDiQrrqlWWsMZm4QTdu/H7fDQMgnuoXwGYZZF
e77dUhQahpg6Uyq9GVozk+LjkDpgzhMNTCsaoaifKy7YWmSPCKCImt70ImvzpDz9
UDe+bzahmQNOJE8yQMeHdoc0pmmDciGySSgthdA1U8TLpesSFn6WvpJZCiFEnCpY
bgsM2KGlPtf8f/3LQk26ackBAPUfmpay+lb2M06vTkXd7VsztU2U7K9f6qUPm5i+
2UUhBY98FNNgxD2Vi2AFxCwmQShz1Zeu3FFYiVsFPSclBC8WZauAaPuTJp+zheII
T49Ue2Vx+lgYXWBiQ8hIDCPyhrr9qMgeztHogEFWJ3pfZ+2ksUsVCKZLZUa2ZSTK
TqttyYLiekjm466aG3Yh2NQH7m9XKbHKm/0o80c7OiNgdXGy0mVfzGI7kkbUrp+B
/KXcLK09PJBwKQulNI5mZ6ysiRohMFiMbizgm2HKEu7yd89a5Njh9iCRSrbMFBWU
oTiHu5WL63XyNoVMEltvLWxv+HdSBZc5uXoHqRFRkZZLarrYbtIEBMIyyVe2+fId
JN4wg6o7YWY2JN92sKlwUCn3uBgcyM8lCjbttTrhOF1Ii7/3sg7jfUtJEANJpDJD
IHiDoLdTW0LRhhwL8Dpz43O74NxRERMqn6eSGe9fhBTjNMXe9aTM9DkjgwO7ffqG
kw4AvIdLT03ezH3emCEqhw9BOPSk463pvIjnqwPNqWN3SKg5Jp0NLPGwT1+t8PW5
WvG2p2eJNv8CmGbLjqc8xQWaL69Un3EzXcJjAnUh+PS3FpBZX/+kV2Xz5NSkxppb
TkFS19Poz0Q+qPdQoMEfhLtqjOE+8y8U2wN/tnU5ocstLUjwkI3vVaXmpAurKE3I
SGhGO24LDid/Bz98KMjPvVkxf1oAf/NO5yf4dwsbmTf1+Icf2oV5vJ6SxsJc1VZJ
q8fpq8Lwi+6bQJn2kR7wfZhqkETisvbXBNQqQeMwIH+HKJWsY4yk+Yz/+jQHX70H
BQvMVt163WCwkYz1Nih+jtnkjA+HNxXRejQcXvTE1x+y5v3PWHTPrj1DnclSj9dJ
PtgfjVekdf2Q+WvRWjtOAQPYPlyafUsvjSJ3NML/sobnGGIJbTlIrb6f7i6Oabt8
GZvI9TNBXEKJyjS7rllC5pNCaMJjG+QamxEThKUE4Yl8oKb4Ud/2J/3r8xff5I2M
SYNhKzusPEPWlM8aW6hC3oNUqo0/216XwCTvqQ9WQToSi25bUZ1wR4EHDQzFqOec
d3OY0VZ1KII8ORLkFbG+q8KF094plPjn02XAnqVrLIeRAHoZbh0r4JGAEOviloZM
7OIFzC8bJCtIYQq4B9hrdffpeRmbfwJFUk0G/SoLniXXYWRSE+rfzx95J30ft2w8
TcsdK2i43ge5QAaYInpuC+PIVcyk/d06HYzFzdkivK1Ode6Ksk6tfEOq9WV9Y5oK
mSxjsNpKSCDtV00R8u7c2n5tONfo8qGJWng51w8NkYSiMWwmq1gYecrOjuSwGnW7
XPhXh614ROwH7C3r1LaY82Z9z7mNaEphlpF32O0XNVabIcUEwc/dYj9QUpngHbjW
Ypq0vSMvWFTrM6y7SmldVjr7kSqCgA92eiSmT+nU01tIuUFYPCaxb67wEAQ3udlD
MdM42Uib7eoLC+ap/nl+TrtMYnGMiXjKjlTzCryzPb1S1GhWlNA+nRx9DyFIxtJu
JZpP9zmmA4U5Fm1pfElSLz93GnAMvdeC15OmSB34oAsoZSdboeu2g8oPfcWXaTcd
4oU577TAr05UUMM4Sz7w+FeZd+7RkGCUX7RdXycXpY4zpjgHwj4u8WqHHTf3l+yl
kI2E6O426BTy/Qdb09m7B6I/k7K9N2eeL2dthW5dHWurQxYEwNJsHOmXwbeoePYk
3L939yEp8OZhBroOcJ3zdKFvAlOsxlK/vsZ2peE+KmHGjS+JAY+PrupkmkZLqo9E
9kEtHtLT9Gl+lgR07Osczak78quVaARwdTA+rwRLJ/yc7tlDxmmjBEXBmpn1yAmA
lrVkdplApKEhd0uMYtgfBfyDP9IoA+9t5zil0d/qgzo9hYnYcLnS2X+gmk3nvZQL
PEPX3o/7J4ZyebaC39X1iLNkmes0FbAxnBxoqWt7MDZVN8jT34RFxVjsWd9t9oYh
u0SsTLWoKCGR5S5yU/VmEKvMOm8wPAP7IMEuXGEiSV1/Gti+VCchpwRcGtmq3URv
acVgNFj4ab+m0poH6bBF7jnx3i+3XjdfAPwGXroX+mck7XYS/qWPxa4DN/g1DRf5
I3VAtW+ExKvxVuRm4IG104zZoAKwkGxcYC5Lz0PSWlQIN9f77OkHTHZVYmoO+k7+
/7y6MBtSuCPlRXdcotyEwoySeyV4FZkj5lRzwczt2lXaCw8uuqWb+yXs49vFU9tE
cqBqmf+5sggYSAil6091XAmM+S6f9YQnZfvUclVI9X/uTmEDMyN3pcP8eBAAG6EU
9lnkvQmfVEH/AoyPNRHmkpDGoXalliX53+ZYt3tcK+yJbuQq1dWa14yI1EngMbqX
Q8vylIiGbmw4kx2MlGlFtkHMx7UZZ0uefbuHxTUaY4L0nuJLpudcRUuoMIx+nMsO
x18kw1iNnR3FjFmksR4XfwVMCAg9sqkacKSRYGlhrtNykcg5ZjnuqhP7jG+okumz
vczmUviOBwyO8dX9GNDSsdfgt0JGKJ/i9DdBVHvgL1HbE20NlkEoDaB35mm2S/M/
EQ8YW4bc8cR3XC1QNvG54X95ENdaCz9N3BnorbUzSAbBTeQCaXoaO+F7dhXW+DE8
s2+edI7QIWDP1vlDhzNnCSc/W1T3aqWGyYiA+7JBY+ynZ/XkdtNGhC9ctqaNSaHF
i0EPdP2BcbrC4BqNuFkwJpqIMIuEEST/s1ajvXkVc/6SAjP9WcpM/e04yCvp0b2a
0lg8luQDTD+dYmNrxRgtKyI/x7lQG1flcXbkdga8BzUubgg7n0e9cILUxJcWCD8N
fa8E1Lga9quK0G8QoaQx3+BPJEowYN5QNjPBjqSbW2ZJPruGK2AiE9QhxgpSUFk1
UmMsKK7fGNLLb1Y9Q1rWE4fXJT1Pn8tfZeitFfmVKInnuR8OCr8UMP1QDS9fBU7G
Z2GiEG8SKCpq5b1TJIi0W3FnS7HNqk9A3TIJa6lfJT5yxP3cu2eSfa2CIugAOCWk
eyL/RzqCoCl/472YPRIROl4fsBdJm/q6St2x7RFvjKR40mDVuIRLwMYqbhQXwSvr
7c5V6vblL1/3CTvumFfqYjwVg28MBiPLWK4PElip+WqMeGMgMVASIinS8/T21AcI
McNVf+1rv9DwrD5cLZ+rSpsjtYX7ej8COpHXLxj+tQMJwRfPpRoJFslJfqjCW0ke
XVMLIC/2qFTVC6OaghHYjDs+UiiPC5g1P/G9CtueLbE7CMOWMDHMuNr3DbdkmlDd
ShpijdI52SWC1eJHoPy9sSEoSZU8HxU2uo/fe7VilvqHvC5flT0+rpIQmdgbPqQb
HCuKvk3Utdf8KFmWMIODoMjjxElp+2piyCYrU8fMfE6KnBPNP1beCByMu5pkJAg9
MoVs3XKKGxqLTLsPjwMolc3lg4Dk53u7U0WUInEZZ4wH3WKcAECDeanptmmnJQm1
n+i0d6/u95f2w1RKV66FFhc5QCdARKBkcd+zDIXwXzxMqS8oj1HpBYDZRPJkA4qO
nt3h3cqF0mmRSUyB8eBbK0kM7aXLi/nBa8m3Pn8F3oKQHBg4PmsFM5XrFCW1Zj9M
3ygrqmEIIqo/wTwM9MyD41RrB2HP4NWOtCw65odvkpvZFIz9N4GecPpviGcOOqM0
NXl1OsUL8YbsMB/1zUWN4aZkFvOexzu3Ma/AOfASghf2mzBhTB/ldn81+gObUHGs
HaMretKC6/W7kKUIlCefdJ3nxjlg+FcawqaL3s58oFVKaSyocsAQnoSG6TnnslzA
6fgCGlf2QL2nRbWYYg231UdswcSl4e6RsGM+XVvxd8wproQMBcImBk0+Dehia1fV
51L21kQVHgaBIe8VaeBYD1HUyPPlmVE9dU8pROQGpOfAKh8CecDXWkYxtcwj2Tvh
mrLxxujPkM5xHUv/l/AGyEGUSsd8Cs52xA1sb4owirJjXD7AsX5UbecM+jemqN4N
cnymE3vJX1afh8C4gf1nHFz67eBNJY9gvMzBtYJVNZ55W30H1bJToBupUgskTB+H
2H+vNfniMyZm21571R6h3z5bcTxOw7Wsd13Jo8JRB3K7OsLqgU1KR68DJmQbBCg1
WWZigtkJ+ZOAXKM1nYmpcyAEBYlP4pK5iuZo8HrdsZLlWBgME7g1GC/QyIMHOoAf
hNBw7aKrdguMP8kbRheXjSaIPi27GyG+n2oghX2Yo9GiSXP8OHj7DWET6MMh4PUp
M4Hq/NPK8isK9987qHTUkJx7+VPMGqxd6XC13w5kBevm7ua4SCbzSy5xSzx4ymRk
RaSGWmlKqL+VYQNO5Rdn8ChBYd7QiS3qkELgc65e+B/HgZgE9EZhDSY/AvDHqB8r
Po81VkTzj6jG5xwsrIUM0wnDEZEI+gVyF3+JgxOfb97SXh1RvZGbCH960+JPIHp6
iblzlapVhu2hKOdm8oaMzLxKCS5s//yQtBVRlWaIi1W6x1w+bUc/hda4yyO2yB7K
YrQ1xuR0PgUSbYLZT0/LJse01cUXN2Jqcu/b38IxJ7J6OJwuuLBsKFgX/JqZ099/
EM7r590/1ly2aZVgEsNnOc46L4ykxbeAon/fViJiPip55g2jyMeNlUzlQlMY46WD
h6lY4qUfTRElCCLZNSYhV5tw2grvvne3lZNEgTaC6aVbaubjTL2rvwLO0UZh1pAm
BNGkRR+of7V8pHVsXYWmt1XFEUwlJy1PoBIAuUzbYL8UUX0K1Pz60SlAKpCCwKKB
sYoQ0uYwkRv7OTsvBUv2U65un9uc2wlpwPFvObOqONyAYy8R1rITTnlfB6XfTcMy
GgkRMNB2yLOHRXx6Jn/Z3WUnU/7uyILd7Nv+xKKI71R3xRjb1foISg6CWyTgCjvF
i76OWvawedPwwGlwkjWe+rwJTf/gNcA5jIkqPMTBCxnpo8/Up24unHXh39B/SRbS
qjuKSFG+y1qLjujKevUMuS1dz9yTPAiJpwEb8KKPNbk4rvwpwAkx1Gq3u/5LGkx0
N1w9cG9VQhocCcJFkHjIGqY/ww3YrybmP+gCIzlKum6r6Djg//BtQA934rUKNN2c
CtB2CCNKuUfaZ5s7tiO/1jX1yd1/os7oqbdrbvxM4ORYQ+47/CZqL8s+z8Kp9Tf2
Msv4XRYdpjQget6VIgjKfdrc/QWuOC2/DDWdI+6hity+JBxbXxVs0R+KABVEbHvf
2gFs790w3T4jWkOHnqsHnnVLoId09yb/UzgOC5ygzoEPRscbiVYZuCibdP+sv2fZ
v5znBiO5Ey7R1bcrDniYwlLm1/+Kn1BZHEa7Dy5vfEbbC/MrPI6W5/Wa8MEFFxSl
A97lTUBadrgjNDyMmS156whDIBzoil1C0BFaCR/qfSuANzo0z3naohkVRQtjuKrw
qE9qV2F/xP9aq7PYTTp5y7fnD6yZPWiUZi61Jh0AH2f0teTUJkPYzeyOJGcFWt8u
AwOM0lEbi3NUZvTD+x2ksoDMaFICTUzM0CKNz0Za9aR08z30yIOZI6vvUa/PFi9d
UAzOZTcDXZV2mldlOhXLI6WjKO2QPgNxOczl2SLTE7N4GxnmW6zdG1Bc7sXf/amE
GDq/ioSlrop7s95TKKJQoyBgMtZZGxV4luCKjCnzJcf/ersdXOc/tw7ex/7oy+qg
Lqz7MbuXFNS303Fze2YHv2ggLk2fFRj3AHhOddghb0Yk+Y6ByoSojK/6Y6OqPo+A
TO0CuUsnloeDIGbYIu9pwWdTOVrKCE0ghtwzhjPANRxWYx1ZhUItQAfWQj3TO2Bq
ltOFPGUQtzYeDIOPjbjOqDiWDh9ergL1hDvUmJFQ3P1VKK/VzdVrDgK8q5riLZDZ
GfUsR4fclWX1DbAIhGjUYgVhUlsXUgGm54O8u1x1la4sPy/MTDYbtxa5gp/44Be7
qSV2hfDhHZZt7UEDk6kKwRlq4cS45R1DM4peKto76pyg5aetKukMYgi1kJC1JJyP
j4ba9luU9TYay1m0ca0ZdcGHJPX4QAHDZs4dIY72BaGKXcIBxtG+x7BP+JpmkYs9
kSs40XanpiB6CJGaQfX+gFKsXb9306KWAHMGIwwyhTYYA0ZHLuDJi9vJKy6GcHv9
Q4wG/sizaX6bMiqabqsh0zNTlgZJgarNRxIx48Uw+LoI2rXFHr7DPsUWuJV6oQEZ
Y4FenMeu+8G1ooeuO3O6JcxpjGv8IXIEy8L38SXXtf2qGFVnAON3IlKoljDxid+w
jTSBvja7z4Oz+OKX3t00ng0Z4zF3X+0ki8UkyFTeNrWhtouIxJomAfnNOg67in3I
GNAq984lI0rN+uDtBXxR7HPSWHX0slQWVJVl3J+3F0TrJYyVVkdhaZYcoHNOvcjA
ef8INJpKRoug54eGPFs4Pj3wygf3jdt9NtDkroXpn8jdeIVt0tPYgLYHbdSyvHJL
4me0di7444GPgtuyzz2uJVv9V99F+R9s5WldIJqYX+aUvNoWuZOrVhn8U+P92wZi
4pfg0qi8DceICURWcjcM6bLbMqdybSVRZ5wvrw3fFDrOnv9qZHOzDpElBOF8yuxK
0PZ2TudKg+ZDvEu/tMPRJPOO8qt5hwD/ufP3i8vLdgrYNPpxC3edR6T/5C2CwKaB
bhxxpzhuNckgPc7SnU6b7vR6U0fP5xi4qZFhWRz1FJe09cKW0e/bBI7BhVYMI0Lz
zLWoT3zauKvkaeeG9VI1Wv6p3O4FhgTOScchb8l6tcifgJvC/FcS6B86Ztg71Ids
KabbZP4TRUXNrDFW0zZeoPLt1etjeluac4pQRkyc7uKqLj82ObNDl7M+3JlNFVxO
cg8H7yjtrDqfV/buynIaZdJQ6zZ5zuvu5CCJh3L0u9cvbS4VElbEbZFqg6bzfI4Z
5EF6KBiqxZYXskCNLrmMdDp2VMcDANJO6Eqt4FWiM3lEnZLQS9DEtLohWhSGies1
7+7YXlljgzgSiRcP+SsP1SIDtUGbV+id+9n03EllfmJo67k5pnOxsZJrcPkQBDZF
VtKByrysbQ0lC3HZY1Cd9Uuo2PX+nb7IWFwgzMLqhlTVl1IzymWkYmV8YAT6XBB3
ZjGPOPb1N368d5cBVIgRHJqPO7ikSar/zmdk+gyYAfjWMj4Kae56T8wCOTKNoF0L
sSOGcnRwYSpj10csReHyO6igD5J4J2DvJrYDXahInuSphnd+SpOj8jwLuqDTpBJU
UTs7IcXMF2BQB4t4/OpJJN7CG0t0U7q6X4PdcSHeyF9KGZgyH7viq31h1aYNjzxP
pa7sQRXdY1A0r05+pIwqcGKIZzBATmNNs1kMVgPXhsc/xEPtQQWWvrygnQOVsZn6
KtQwe4lNyqntHqAsGhW4SIj41btRMwsKP21vjlU5NHWvftak3PBQ4IoYO6RsIbQA
+KV7HMCPKajKaC/ldKLml5KWB7u5B4UtDgo+BIvh/LH9lef0tvK5mnR57+UcoJRy
k/iQQapWpC0TU5+mFFooaxX2h4pl4AbVYL1gRKnbXKNHmxaM5piMd/RjaA+mW5bI
J/z1BG8sXV/JNcUKO8OyDKyfgqp+slpRKrCimH0k8FtgiRGOeGUaovI/TUbVk+pl
lFjY28qPNho5H/tTpKkOD0od6gPCjxWMu97O2QPaqZgsebaOh9IkbA+5GKNdHru+
K0v538JqtqL9kTqnwyiCldVvKqT8XOYmj0AdIGVB6zHYz8Ntkv/ECYRXBl+QVDmt
1XmGWvSz+PykKDXcqWosQDEUKyh4oCHUsRL4X2CzBLfk3zxnc6fDV60YqNQ7s6Rc
dB8N8+WP5wlDwTcQslEVVT1zwAi+7BJxUx8k1WvldnGUOxo14OMs2eDnpD+jvip0
EP+BJZu0cmKy4qB8Joj90QjS5JYzqOI0oCjMrNIvoHzxOZxmhsddm4vfmi3ZRFjn
fqNYqfRo6ZmavfRleNZuDx/GD2Pz6d/CxFehXY2tqIyRZRW72DYuO0y043eve2jY
w0FzeAoMb+PYOaD/n06sD6x1yELCMJqaNdqht8mKJaXMnm9U7n4tSErlfbSrQVxZ
idF6/W1NBtHX3xd1xSljhERxZKLaBnvkKeW6+a8jAzhNR3+YYxhaAk02SCjsmEbm
oO76qrE9M/oDvii09IhLdp1AQrI/HfxP1EhM/6x4PT5H4vfnInWhEHsmzNEJTsQ2
c3i595FyitGqC9/aUDh8S4+0niSBtoq1ptY/cfVO4sFQ7S3ogovX2+dcLaou0gHE
sXeQqdyRPP1DrJLrnuyWI6UdQ6n1Y5yKcV99IH3O8EzQ8Koh79vbvLv8vEoxnyih
ELV8YwkOYa8DJyCUFQkUQKk3uwJwFaPlJbIQriGrBT3TtFlF2NOwdzlyPGuSOZeR
R4PmkoWCeU66Qnnvhk+sYAHL1AfdUjzN3QvGIBbwRkSt4v5PzX4yxZryi6ptiskb
aY+UQicRpCJalWhQCIxBlXiAcqz7AcQN5EPHqgSW3NjhmkK1r8Mrej/mTJj416Ql
WBp53/+h5fQgJFsDapQmyZjwcU4FG0nM8Qc7csDJk7XTzrQefW15Qz6ECN2O40Pi
786xfNoM/TYgZy9/SLc+jQ39mVGqKBpyXofv1ivCNLJmzW80ypnT7GrqQ54hG8I3
LQOwaKBzBRNzTmzKA1JR3D3hx+XbH3m5OjMa8QnDtYZoFIxNFULWsBlusJSi6CZr
p2leQIORbAvc5eF4DWiQPHUy6FWwnVXAxEzeWGX01DtXWEqo/ledJnpQLJrEyAxy
ffup4cziXQBrRngJrRf3+5vlgQH8uzcHVTmsTEhq8jMbMPM3Tdy6PMjoYe9FQYR3
JymDRyA00dIakFR2p6tciNqc3ad+kmdxMDb4M5JK1jJPqszvZjWy+a8gs4LX+8WZ
qAoLBu6MlpKO8njqSwSDBRhM8fYhEB3y590z02oXG/zSppZVbhpDf8R5ReYlRCxn
Su6wDtXTGG6uuVgIq6KWmtuIXIkSVDHXkqxBg8H1xHXSDy7j653cZNGqSvbgaqxw
hMfoN8JcyHp+aDObF07tz4HMOK2Uy8o4Pc05Z5dEV6CWsvwDYOCYgh3uXgbvSdSI
pIgxIHuyqMKPiP4z+XrKZsZjf4uiPBDuyhHHXo5JxXo+s0NEuWM6LNk8SNZAUyb0
dKHxbM7zui9Vlr4LjHd/40NhEyV2Q3myBjvgme2KgPgss2bwwMgOnD3BunCi2QdD
ZQ/XghYqPd6+2sP9udC7VhBLykXOcPg8J+iibAmhLygdXYunCNxYFxRgpU9+FuGH
DkEpxlwuQ32sm0HtudTOZOWGBPsDulqafEkTQn112NrBVNjyyWSE7jgEXaRHYeF7
NNvkcqETh6eKBd2yOdVlar2wud3or6PO6+k5j4KPip62V3chdaJOOuvi+OuSrtgs
7QU+eR5S/fLemOp++aPgR+CDoYgMcNfVU+EgNQ4ZEPN1pTg9OmH8yUsTTH/yXYrh
pln8FzeiynfarzCjVEx4lIJeT4qkCKu5PqxpMrDIXnh/XVqtZI2yggqgfvs74vCW
hM65lwYjo+WTeq6ndK9ANSlP5beEKPaUUHNInn9GjJWcBX+5ANSlwYFpQmuxXTRX
VGeZy8xdYQxvGSmSch+fpR/+lLfp4bgxviY+LuotSe/kJE7lqqSWtFGJdtDqOpQS
BqcK6Amsk1jP7pOQzr1LnyYGnKiRTAkgiKVDB3PKdVdkkCYGE679drbJRvGtWhJL
hA+UWxxpkHr9jfEkC6wfRzdGpwisBzb0ksuGcxJw7yNBkfmAVls5erFZVQ2GIdJL
IsNHqwevm3SLV6hld4vykunV32O5a+q8q5XJYCHcbPjL+XuTTOOy6baxvEKOvx+8
8lP/SuRgQi8wKgnSrciZY3n1aetgeJtLMg192zPRTBkI8FTyZONvXO/PrJyyEl9Y
R4JTFuRDzzaONHz553LOmpBmS3EZ5BO8CN3v7bKPhd20uzuEVkkNry1pC/uenq9O
y0z+/gpQ6SN+6u9k/fPjEY2dmQfV1f6+Ga7P+5O9aoEfdM9xDptkiaFSBYxbdY4h
71pP4ehiyAvjJ7m1ayKxtQBgTDrgdzPN1oGdivkHxdWL/D53uz2I3rlKTn620gTD
EgXCMFDY6RdGwDE9xZC1Dn0ds1Og+JhwY8NvR4olbC2OJkIEhRqcq/eXYBipk5aG
sfEYp0DLHrRPO8ldgcMJ1BAme8Z9+VhFaZeq8tUrPHVhfH2TZ7jvGxdLw30mMkhq
mC0jHIhILwXqXt/I2xw3nfD0DOCAM4mGgpKizEC6l9L1z6GqNreIl2F/Mf988NYF
0oBOIgvR2hKETNEay8bbIkj0KyKDl92Dob+TpPD1TnknFSgEZckiPFtcR4ae4Yza
zoLtejCo8GExv8zbLfR5UnOTsEbdaMdYvhNEjA7jKUc+1vUxcma0OenjkuOSgUkh
5D0lKK/JLozOZQiW++WxRq1IwsA5AdQep/InLXaP8ejhTaLdnAmQLynhdzdYWeUx
WipYqw8khMk6Nz/mTIEuiBIWdYachj6XXUboZJTWeFKaz2BJ8JY9Ju0rBuvT9w4B
g3lTQemcE5J4WxjIIJhLaLe62RP7LiwZcLyKPKLHvlNCe/jHnPTufl4qeGY0XHfi
+BUf7pF2xGulCl3TSzh/kBabNYCiVmx2M1Q43ROYf61L6M6KpMCQ6KQV9BtF+VqE
JRbdYpvmM4WpeNmFpma5b8APjybFpEp5TLJwg5wTEOjKLKgzLIDAj2X/zcHzgmmq
MjeKQnImjNYfoFh070CNl7TZQQk5vss5oZK+iFI5gkjEzJCy3ePTtQpV+m88gk4k
3JEluol0Y1jkwGz+X3oo2ZK3Vmg2DwcLE9qwrOZRC5GJBUYaghxW1V9AHKNSDjeM
igvOGwnd2IkIzS9JhT8l5JO/s/276KORPWAxagWHIpbp6Zc2RgseoJ2xkIMPNkec
srCdROnyQ1MiWiFVueXT9oCi9AgkVpW0n0forDJJYycak7ifCrjay0Y88njx0BS6
czeBnbBKBCPkVxPr6caAIK+8eFVjWaXRvJyKpfkRr3KYt+QBetYjmgl63ZiNgbds
UdOPtTr/hL33+rWYmKKzWBqHaWjmDjuYlbbM35UQs2aC3KPy7pv3s99cfHK6yNlh
TjWOQdm3eUcnu17CPWakDmlcVE0XpIuVWddpYRgAbd4MsMSHji8TpPvCb3GzltzR
TBl2h0y3tU6U5UocdivB/v0gCN/wG5ll1xJ4ollSnlkr72dgbPOZ3B1noo5gl5/O
YdYhP5yFU0b703gd9HKrEBAXbG4S1A0qVB9aXD/WENESymRNHpXE6r8O/sfTpUir
RcJNfvIBwqlcgeSZTG/9TeOSZel/wEZmGITBPD+0552EHAgrYCdHA1crYdURJQqZ
4XKoyyCiYjjTjxEeB7b4lu34FTm80dTYzo3JDRQjamxWt/8+4mQa0JL9HeUK4G9b
ycOemnG8+BTywafCThyX4DrrfFupR8BKAcyBD6VjLmr7BmxF9dMBKgLZfZ7e3XVE
Ev+Eiuca6HN6UUuHgsHMAHh60ZsUjDwGVN8Yd/iOJ+jodydBnYU+trBLr6FYfP3M
pQTUOM8PPET9moaOENI+mM94IpVycDKyn2jDf3PRjGGdFzl1swIVFW1D9VzhpC0A
vU1DM4KC8ohHwGnGZjmaxoJSxRJ0rUVA9bpVNC6r8e4GQUaobUc9SqMLXxGUM83H
a5LItydj9Iyr0uD/xTa+DFzoFY+DnVOHmTFu1oPO7E0lsVNSffU4al3nvDpo2vze
wIYDjxbYW6howm8e5g/q1D2z2rstd37h3lIrucm2Iq1FWlWACdzJAtpc8ZcrF7bF
h2H2m9wbVFSCvBvLE3DKpOXiPAj564ms4kWht0foxYjpImrBMJ24Vi+1eSFn4u1r
fIb80/NPROAOQMQ3/LNEZ8Wy25lfwXbSHejZ54o2Chdyofhqh1btiolhjj8GoERj
198xDexwr6llPjtXMHef6XKfOL8KNBXz4be7MzU/tWR+RovhhHpsp5iI4lO3Sz7w
prU/mOF20V380x4JVWqomsdHZnJVmCh6rzvatDia/t428Co6K9mr7LSt93nuIXyX
RoXI2vPHZ89O01EGkoTOc0S13r2wzADL2sRpEuFZWsbXiSggPanqkMspJtD9CuXN
iFh8ZNEI/Nkdpb5MjOa/bjXj32qprgwyb7aoNsZYQp5Il6aECaSL66iF3q0STQZB
kENdMGWAEj+19jnWtsFWXNB3LkBOHRvVeqPjsP7khUdpScIbZ9U3ruQ+1lc+PcVY
iaIA/ESTOqEycWWbUpeJpeM6Vn0ykc6+ZnQ9evYRL5WSl9GiSqucTtNdw5AROcb9
VFt5KmmFpyjyJ17P4uoACKVlL1K7SRNTrkKLGubUEPlv5rscHTAUCbXzH4EtPhOf
qqRvyXSxeuL3A0nm6jIL5mfuh+rU6FDnCMAvsxzdGwtZ/grd3tGca+NRpPBjdNJK
avrUsrQOoEJkdkIR17UyT/dAdOLvj8MhT+YocMPe+lfE1iez+/LK+YrqHYxh6h1y
kEmZiDOjjWnmJqmZXe19zsxwGhODu5ayEk0i/HKrdMA2e7/c79Vv9v1ep1ye+hUu
MSlv4dCBgpTRy0jbm3ezTHbB5tdgVkHsITrnWACUsJPju17qDvt31Lbs0YnfUnG/
0NphNpTtOionw0NHsD3UgcKTBwWY8KEsl4HehJ8H/4zLJqDyg81a3a6BGZJWh3/W
bxWeow4piiKryb3OBfbDHp3IR2EITr06eBKDeileatVuZuzw321OKi616hxPkp/Y
qWT8RIMRDY8QNetlTxg0/eW2UXJgwU8X5NMAq8Vw9JmKEOlGgA8l3Fspz+iI+y6f
+KeYsdKp40zcSTWbzJZ2hn96xpBVG5pozLMMPnS7zzLBPo2pSYo+ca8tY+AFZYUq
bdDCK0xdec0c8KCYnNP4ndf44Nu0T1xtfmxDnpVmP5W/+gBV9f3Iqfeio3IU+ZIF
lG4CYSA3mv099UXIsLXARKbxoLQi+AdWMWFHnS1VCZG4Jdkc81H2osZ2Go23bZJ2
/jjh9lPAnAgiwWWDsZ65Cuq5OiNzKp9FgRlLvz7xZRtjbjhxC9Pm0xQjnbUEOKNZ
d9af5hfXVsFitOK73RHINiEgVr1VMlGurpnBce3FP06e5cvego9w+ugSzUS1piLa
YuSKVjC5wnyNsBlCEBJJtMdhqpkGVPXCprsCTykc6zhGwSK2nsK2RIAgd+5RECXT
zLz1uCDGGno3psAZ/DBlZAK8O8f64ceCPim47iAUmeB+XEsQGmDZeEspCwR86OiB
+9ppwmL18pmBNlFyaz1hgQGcUXLR4Syfmzu1JDjNizqnKAU3e5MMoJumYyOZziHu
V/cFB5+NjbKmPXj+KrqxlUaWDC8f4uLH27PlD5sDR4JBaZBsKv2/B5uxyD1Ijlzo
RWUi9J1J4lH2Z4MAQmyecXU4/itHc1oJwCUZjaajhOXqz6jOLqjkxu4BCu1Jvdtz
ClHyCnD97YFeKfwe36GdsEp40Qcb0B7BGl4oCPXTqOpnB8Ohro7yr3vFW6EiS3hG
aBaOjmdysX8crnTuE0WuGKJ4PUf9xVGbRWkKYlTm80WULoECmbaKRuvoiL4C/skn
Q9BuRSfglsZp1tY8cOJB6/sEfOl6sVvapF6xepM7lVBHngtA60rK9DyEY3advdmb
xRmJNzEo0/ZUoApYwjq14tXIsI87L5zyUds4KzGgAUciimWLAYy3MpT6hhRT0Vmr
NUkpKmg9Wx1bLVNMyHET0NnVvj+J5RG4gJADEC6PN6Sfb3CvtmlVZe3igBQALU5t
SRjQZ78yDih2ZbtEuCB/TIMtGG9O7c+ZKeACcLouHa/ZHLlLnJVBv4ejUE72l7jm
stzbJ7U+S/8rdVCQd3GSLCfjFJjQMkIQYnXmc6rAUtGq0lRDU+Mh/PFX8e04H1R5
Pa7YKg187XMN1eMtwQSROfJuGcWFN0MEQFwKUKb+bzJDj3kKoCqEwPOXkGN6hifn
DkQOZuFz1pD4RgWMQgeNIOzKK9NP4YZAuJhZLzqoB/NNpS+orSswTFOcuYMAGvSy
Y/Fvu0J2AKwDrkLB0wBQ3zDoGCz/4DtKjtLMxQWSjxEIHRAaIxs66Hd+sWsRwNVh
lTqpLEDiRg6NJKAkbOlB2AGcY2LbVj/ZTIzrCsW0PHi2dlQweehg6B+R5kFZ6cY4
GlRHPrhWaePWpCg9Ssx+ktld5ONRwP11HtF2muH0Jr9SUIX6RMxVXCQYJe1+sT91
3QCWkFQr0+TSZvQYmg6E8ozhlerpwd0pBZOqKCDBK11Qsr1inw54KJYoKlFmj2CQ
XwBlBjNf+aXRMfSQHXbbY6r0Lbe5nRexsQirW+KrlEJVzTvdupLg5islYrSl0KwK
Vp/DF8x07lQaqwZdhUc48gmqipJWxQU9g1/hokmOkO7pJDYAxRqFKQR/XtE/SWEu
VoOwcVxIq0KXqqbW7v0NF0P6iqTHXbw6heAxydvz1tkzjWcdSGuyOw/hM6EMUz2H
nM5GJ0FchxeXe/dC7B/SZNmTh+YYlFyMjD7g9Ar6iO5pZO14/oV1jOQAoTtbN++q
rokHmYblyjxlslcqaV7jtAw/spYpyXUoAbPoIp/7yqkTWvMG99HwWq3Wh91F5GYp
iG4gxZMFaIrx0O6LtK/P9V9hjdYiCkvVDhOHjTSAIXf0hM2q6H78IV6cZyUzXYQ+
lWnsM9hoPiHRVpaRLMs+wStlYg7qqOPqauRmCytqPg5z0usxyJJHiF3eLCj0vQ+I
LGjeGbHMPXJGBJS+FirqE+N4NX2otLPghgWFDz/oMAu2nKIHVy4N1eNZk93K6CLO
qNU7M4512Jd7glTzf0wjZ7sbJ/zS+TEsXxhmMfNtqQzKeV9q9Nrfy0VGvzDDJFt+
eBFV204/GZd+V6xrzjVJatN49O1KapuWKl3CklbFRzEdvtmMbRlzSVenE5Fo/GUD
0MNizCEf8iS+PhW8oCBfepMc71mxGPS81VFuR4GKzNg9UfFyFqZtxRTg14EeE5ip
Nyg/x9LOk1/Sawf+NqscOromeVU5Mc11aN0I9NAS4VeNxCF7N7qfV1lywXxSooc4
ZTFLxvUN2rPfy26v0DoLnj+fyvkeyAuIP7u41dSt7yzl1t9jAPPfvaryzpUvlh/z
8nQ5Y3wPzZG5bWAcwzgV0/hqAedAh3V6l+ZsCQEmr9yKttEeWs1KHlZkFaKvkZ1V
3JyxjWcdga/SSfwqo9VZ7JOeQv0ICNZVD+U9Rtgvh9e+zQR8w8xfSIFeTZ4DtzbA
DaGQToLeY+L2Is5QEaz91aw5GfWSX/JxzDoAoMiLIiPEKrJR0kCj9ECYjzwuM6bJ
/E+DNGka0CiOAv8FZR+MG8ZssxtxFhm+2n+QxMIeUMj2rd7ZfIsP6sz8D44FKMFy
yvJX5H2u+rWqC6JOMey3/Or9oaApYZ/HyFl+sJWd5InJA0l8MIDdXX/rpGi8HOtE
Ehx7DAooHKgAr44XEtiaIgXtoDX/XWBHPkHaZ0iDIu50uj7VClFcKFWUfUGktiA6
O4Q1AkI2Q5Ws9UBlqS7RMkzJHoaQiesl1oaL02LF7PJN7GOQLzMqz+I2lYS8LMzs
oBBFDZPFIskVYxNGqI9+1tTeaMjcZIgri2DOlARMhb8JOVLNeXUwqRcDsSfArtNU
OuNdiqFK1C20WtUxnZF86xROJyKQgLMlg6S7IzC9BPKGfQZR7WuMLeaNuRI4k/Qe
9yNuPnr57uoUDDbf8Druct1sZ3xyudLlESw1H1xNWAIPE3VC36zVbRDsn0rrqRUJ
+vORuo43I9PkJV0Z46u9KCPBw7pmbm0Vwtoi72941UoNHbkjVhvazovlAlkSg7aD
4q8Dy1abals0ky/w1O7tzpjDh3TyCyL7BoiYwZNcHiaOKXd0BpLiPx8Y+4fxyeeB
oPovzMm8aaNbp9roZVGRdalOq4oKYHJq8pwn37U6BS5xrdAtDo4LwjnCKKPuzDfD
iabH65MVtyxSSe3MLBjPRBuxWZ54sn2HRBrF7ZjbeLBk2YdZnn0bGcbu2Ahuql45
xZ/0DVXqdM4xVqL0jJXD8tuom9+Ep8IX1wtBbEZ42oJBvCujXUo0Ae8byLndAEhn
zBO9mbeffcKK/mG7PFnLm2VE4Oj2H+WSnNxNI62s2PodAXYQyv/drvcBmE3Twp/P
2AEvS/OYuFoaSoYBfMLtw/j1u2cdeoeXJ9oYdfJVpE7b2f9QUg2ZyVllHn7YBJC7
grfD7IeLIuVrTyZ9cfoMpW38DkDCz2N7J2MXs68MHy6ncnNtXeL24zK/VQzORGAn
B/qHe4iKcQFGjj6UzhMSd4vIu+H7e2CxSiB7N7gAYzFxGJNOycW2oT6BAV3qoiQr
x/4iWDtuxYYgn4HUufTFqedgN8UgjGjwZvRkSVlrY/3ELeE64RGYbgTXQq4INa0q
U8XFBYllRa6XmA6gD0wuiZxzQoY265sjKUjWvy+Ze/hzMLe7+VMivoNYBGFCKhKE
abjYJf6jV+msGoJYlZMuAXOkbQpM6TOPb7ijc9Bco41e14LlFQQooxKIS5mKv08u
86ICmuZh/FVshdZjRPivx9nHNHcDOkuF2R4rhfIEjv0b3nJyjcT38vpjJoSftWmF
w+7RvmHy/12+Tnm0eLNKS/DiI9+yv8jmZwR7L12kD3COupYCBRh/iNa4+G3OYlNj
g0gvje1fr5aD8CxoLs0Vsoj1FyJi498wXkASlyGm3OwX24gZFn1L8QCSeURd7P9D
Jro8HxN77HiBTDEm1z3oIhzyetotG/EDtgF0WVqqz6sU/t3WqsB3QO4jYk9U0BQe
istCxM4gOjaRn+OnGe2oiMn1f31UzG80fmTboUpg39bFvTMAQpPZtRhbaORY07gf
ONRGTIE1hOnc+Up7tcaXEh0+DAAO3BLTq0dR81D+I3KCxhXnsodzPckqyVskQXga
eEiZM/9Ycshx9xysLWi2w/HMJyZ9vbkVk7ICSCaMpDF3FZlXg4KQyTwuIln1eMj3
IbHk+nPU9Emlrv9BEWx4tEb/d9u7qpHTVcBYybwpC5GjMmqWq5pPXX5Iu4a/XPxH
AiHTgETGlbX4T053hnzMffW7/t8HNoyfZwEpuMmJH9j2dcc/Xcgp9UiJoNBl9xLu
otSmxzXmQCOHGK9/ki1hg6D0C/1ehVJCt8QQDg7ETdfjG1M/aweEBTV2N1OR+8Sv
qKLJUDWJ1ZpPcLSW7hJ3+8jrvp+ItCPLB9gIXjhaD4al3VMiRKF14pH6XSB3UAnQ
1pPUdDuFW2RYMlqBab9OIOiiUBNVRK0HHDttGN4BphWIdMu/7MnQtAlXTywTQNZC
R+P+xUf4V7i3tUd25J5NN89xhtPoT4AAulu88P2k5QQvNPgPZCYJ4Cc8fgEJXngK
e2jke7Q5Zeedu9DwYKqytFGvBXPrQ9K11cYL4JKQv1QdnjHP5eCPtcsPVBs6aSau
nYS5GxzOwIzHiUZbA7Kz2d8vZccaXz3G1B0jkRQ481RDIFNY+jPGg5pqOcC8zmpR
Y+liZXRrwoOE1s/0QqROxCCz5kd5yT+ynVxr18u3CovqTGiHC0qeekx/zPnZx7pe
r5L4iwy4QNIfOjbXqhPGaRObRwfK/KOwB8jUsyMUCALc83DMA6OV0z6WCnbUToDS
A5wTy7omIkxHSbcqTm+y/VxDwzvFED+ajPbq2C3u8nK1+9HNToDyn4AUANjHWJaK
MEAaQqI9vaEQ9/Od8ll1rJwJ4MAcy9AgJ7VzexE90uaYVpYbUfyB8/sLhVx54Bgv
8qecX3rf4ZPU2mqHqP6pWgXLoQmhtnXWed2L2CQxenTv1F/IZujUWgAgyklm18sl
nejEthLTkwz++OhLvD8Y34Yx+WU6Y1zd4XREh1rpTT77DrymqhfbBCc9lg2IoKPG
FTAyZhZt9n/fBRU/AFmvJxpc5/Pv7zvJraCxjmWMZz91wbkrjPBwIctuWsksf/26
YG4nAyJHNJou9hVNiMJu/qiraYFNU2fB56eM2XrdlHDG/Tg9X7iXHwnVSRptklK/
H09WxiMDF9bdJXJg6gThlXt8NWgWbwJ0A8HQIofkSceMSyRGzZueJLCZX/lo4OjD
kypM7Bq7+BJQn7mE48eil8Z0oWIXwqAMO6k/BA1t8JnyJok2abi1ANPxxS4mQy5S
P/TflJxKO/ZyYa1lz4vJaMeAcn+nxe9PixlQEIzmv8QDln+F4NFZcplhFeQZyub7
IAByEqB4DSmIGeiqRGuCbX3Jf8JODIRrK+A+UOgy8S6oVqCuGYybQWQJTLbet3Mr
cpUz94tetnL4QNRXCZsqqQ3CsXS4IJvAqVTAXIJGfBdNp0ZwM28ntIkBT//6x+WE
VUZb3v4Yf99H/Tn9zVYEbAC+GTlO/pSFA6KN8T6oyJIoVgfd07dYw4hiKIEPYacu
uUikqlr7dD0OrL4EQuTE3oO0Wq0m4aPAsfP20KkwUup6GGipOTMvKqMGPXwXfaXA
rXRXu8hbrYE8XJqOblB35mXDYuboWGqOiIeXC8O6shXfI+SuRS7xKd7tWp4eNpy/
VZ0r5hu29hbPHTPVaUnUSITDebAZYJnzorHsUgUFFiOamj35L/doA8i0brQDe+NG
w0m6Tci44ucktuhRQS/rl2GyZfdR3+TAGHmEzmYXfqxzOywuaVULv8oM5EUZft5J
qW0+iU5Gy5d1X3mHMw+Zg5wPJQSVujgUGnAauCBUqowYydTAHq+8tKNg3OM30ONy
V38b9e2HGaC43xv3cxjqHNKWRtHP4rmrOrZUgNsGGIR0nAfw1Wfh/HOCYGZdzoH0
gxzGjxhZNDy2e/tMvHYYX7Dpr2aEQwyeSS47D9ii5XVlvGfj/wlsgbtQ+VEaflHh
ohjxZlZymACP+23K4SDJMPnHOqUSyG3QGccfWx8pU67bR8fT0viRHHO5V3QVcHwV
zqvNIlodsKiUYADGxsvGEaDcgdzRB2UnzQtRvoMCGMJNI/r5saDPbae9zc3j9IBR
osD4zgjQrvzpCfvvslFRcTqKztg5cPhZktEuamP7iv2+aMreN6+8v+NAvoIqTNZ2
olUZnjebRhAQJC4qAd1PDNODhIK64VEDTu/CLXGzn8lZtJHlG5cGVPY2kW/FLAxN
ipG0mU3NIeYMkpQswY7M9HO0XDcm8o98Jrlkny0u0aCnu6JERHwbZtzvVESAKxU8
fBPHIpi8OUrZ0DcGZ//MwirOk30bVdvAlg8Wuzvp0aOVHVo0L4IJrAMyagUl1IJh
QYoR4IPEDFsi5UXZAqB4oUoFYgil7e/lrwEwP1naZHUzMvvrcZhmS65oYnsCOrjW
1lw+CILWFAZXwRmu9OllD11LCjZDB+ACQsL9VO1ktMXNt9IaXf1j1qmcIRf69xdE
G31tBQiwdJCZ/Bpbrbday/SAf7eMV8K/BL8WaXqISoXq40e/6N9BocLTLwFMXidw
br0kekGnk++fnceGASw9SdHhm3Age8aD2mX0MSf/6XGIa3ETXFp9tIh/PyGbK112
383eMdtXL0z2vaXw1gITcvF+xkWG3Yf+m9vahLc64B88S0qrEZWkhdWpV8AAFUv9
t0tKEmJnySOn8+iJFPTy+HrylOCSNte0G7dkaP2MeidstPTPbW7bneZYlPVRHw6v
hB2H0Uw6cfcPhHWbIQEErUE8NSQj99XHHl/BgXb+L9FCDZH33/FFpqkpMuYBT0FD
RwhTlZDSnNOodQHY2sxuBDuFGdLKMQoJPgFdUUgoDRyrgIIZaByxE508rp9WVSGE
cG7n+mBj344IRYbxZ6aG7KSSo2ZLLNf7afzT/yJOzK+vOtmWzfH7py6hf7s3xKYC
/UQtRssc2D/GSrRfwJNjRfCb6ToULpARKisI1q9q6hkpBhLwTmbdRLj23Y8dO2Ki
OzL9QYMEWm6evu0/sVYVytqkHAEvZeQxgqRXJhkllYOGgwdyi42GKstP6e8gTOlb
7nUCRmMzis2b5B2dYHUbqO1J2TC248zUBJFtK0JARmI94OwNdXlOOLCf+VkgL5K1
wdZcpdjgUlHmtruuLlYlM83Jr64lmLnYUE3xErXfHrnQ9N+zqs0E/TkjjrNpPJCr
U4qBbWbJEnL6JXt11RwkjOTNJqeGT8xZXs/LPW3ChL9K+pKDX3hl2T4JnUAy1EbK
TuW9NLVbuOS20CNhjygDLWKxlh2+YIJP7SuacsGfP2p4zi2WmLQ975khkojTFmjd
wPdD1kAr344DPW1n44ImbYu+FZ8z9jiBlMXcmc/9ejnZ5xaGi8EgRTDe+NzC3gVT
oKUIfV4lEm61l4HOXO7zflRl4zEihKzIP/0gklvp/ivared9a8eEIf+fKJRObRWV
awi8eY+IECch9Z2hW9azMRRecYqpgvgmLGaneCoo946lGDyeosX6sGOsfTKeHBCX
/UvzBgiFkLi4wFMgFpOH2Q4Sc0eCUAbBAmYiO48pcroU4kX4+IwsL8tvp+E8lH/F
/scz+dDzeNxID8KeMwcrWXesA2rQvWqHBGtNMjPk+CfdeL3eyXWiPAaWKimmoX4G
6AdYbXlNXfV6sJau99jvlCgOJpBlHc1PxnsPPNZAh4QUSJ2hsH4ECBZ7pYPW0PXk
gxzV2LJgqTJyIa44dkRqbrapyvZridXy0PggokBIcgx4ouVsETaJXAL2ksAY2L8L
sMWzsmTo6o2QP3JZU1xNzqncs4cY5RlDMrP2wEUPTzWaYkwSBSx5OVEYCSiGsbNm
LUlfCmq/Cp4epc7srQkCO58lblRQBxRod5oIdd7NXeqfzsFv2MIiriFVFENDXEFn
pGNGzIBLgQoZVEA/ALhwA/7gSd6p7tgQgGl1KVjln8AJpsErSE0CzxDQCAMOowBI
zt7uzL9Pft+NtsnPIhkFQ4GouBG9z7XjWh889w1hTEcfZnDTBOM2+spy5KzQVVRv
WOVlz+VuZJzynRce17KZQUvEO2XxPIlJ3s6fOJV78fd5rzctSjAAZlsar4F5AsIn
32J9FAa8KK4v73wgMcAy0ksHy7FdB7YD0YBCqNedEPCmFX2BwzfX5Yu3shqn4M5y
ZQrgYauJjoha+obO0K1MncTVRk/sp371lgUn4QCtWGpOYnR5LplKrEnzkzrYemAL
ULdrLM9B0u5I/gj3EZv0+1eDYJtXP5k+zhAPlk1uTOPdmTQdP8B4IEMzpi1UoOyW
UU1ietS9LdBd/4A6Qg65qg+enz9P5hyj2fFA1P1n1cCehEALu0P2fg6zeZ9EVIAf
tHx4oDZ9rSzP6DbRKIczcpKKRddosWLgyNkTEUkPheUCLM5TrA8+sN2d3zdyVA1m
VG9hW2j8fnxyW3aDANP2NUxrJJRCUDLa4o5M2r7PQHUw0Sy7k4PV3C2+wjS4U4GW
Fcg+cRFZfGHmuOCadDsdz782Mj+evTG+UXcFygrqeCmsXFj8L77199KvQOhKpunM
+by1Yim2F1aZZf29j93A4Xg1O02WWiJNXX95SU6r7UPntgdiF/ZeIhEsFW3ye626
Y4d0CBbxzinqF3Kq6aLY4eNgANzJ847PIW62B+kCIcQ2XOegongB/UWA/9eszu4j
iCHWsrpLCO/31Y63vfLvydFexQ79cvg+zUqQPfNXxMVM4rwvahXmuUoqY6d1EQJl
BkyeQNW1pcFyUeYGxZ3qfSMQB2lEgBg/ri+jXk2q4YJhCYZhl8CvR+ApF0PIzMwi
EU/5LxuyRWPLgwOMf2R6i3LkD4CYRwXJjh88tskzEdE+02l7pfUnWRpu4P7WwmmW
HsiUL4es8OLEuD18inmLoLLo0p7JHEnAKWj8qruHjdklb3t4wkNwhS7TSCx7R+rJ
d11ncioPA0l/waeOIoJZI5eC+KFojzLAqaMG+7pqONuiUkXeMrQiDJ4wM40tu1ja
tq2DQgY1dP1DFrj9Wx7kvmba1ZnoLnfBGOT62CcHs0W8f73Zf/dDiuN+aPNS1RCZ
4Ab2PlAk17OF2GBmA+KUKqLyeq9F1Kh7t/8dIi+xFpRWffEtHPbuClMTXNStSDJZ
hhyA9z3w0HbMU/VSwJON159poCAgZwLV9+ttXd8rsIVrpg4ej4E7Aglhx7P+iZUX
4WqVobFml/3b2z4kvgdMJRxZKreG7lYgXhFmZ5F/9dYY7mlW4303f69F8cxFS62I
uK5xCsakw0+oP6MsaCuKYwsqp4MQMgNTJCkNoBxYHlx3Ic27ZFEPmUWP+KurmgMy
JtYjyyLKsIqTzAvF6uD+zEOitG2K3hG8KkZf/JIhg6N/0ffxoht3kQF9A4s/Cl2l
pCUyz2ZfC+zQ5P0b3Gr1aYDqDCq4iI9ujKGPwx8ScAMVFcmBgMAKubnuUjPB+mT5
jHIH9wpwM8wgvTwaUn2AuJDB8ImpB8hyfNCoKdyUasGdvoGxOwjrRuyDdEo7JyWf
f0nxypIjAMTtwcJjkHCikX+kBXdkE1Ed2+T0pBuzzBn4OmCSl+sqc8dqSbWzw8A4
Tm3GFVKd4kjemDdfAyuthxuTv/A5dPRuyANXOSWkVaxbL++gG90kpSk71HGhXXZv
2fqFiFnQuqe7p1DyJFF5HPRXg8zD9U3jg2wP/RREM+M0W/UdYgzMCqrO4jwrpFku
VXFUgRTIQ7PZvgDNITkUUogfF6fo9rvEOIcLHZDiLaVWfyH166me/h7zffKwaFth
GCmC52JcWNippsM1vcf9YcFy6jRAnSfGoZdm/pPyeKstCa9LdigtU+ge50LdS97C
gqtSMWF2MVhhkLyLrQvx/edSyA3XP4rg9wHKgMAR/oe6eJW916qxuRWn6axbtLq8
7dgU6IQxebn+/POISngc6uazkzQjwAPT55yzEiuah8HsxLf2+4mMarFTjL2rasv/
pzXJgtNXeO3rVKi7cA1SDQp46+RHWT7qrd3fD5o7yb3+Yl+xAwFRZdtp7kWV7Hvq
wwWUrdao5q2tfIMTsK7Qy/L6KEiJ0t5LLq4u1mEo0oo8NRlLWii3oAPXPG3j3p2W
yldTDdYxD6N9yPC9XhIxR7WV2IWEKZdWpALebQFlqo37hqgWbO5AgMOb4FPf7rW3
Vi/wAoFHRzq1c04iYOieY3wMbxQsEykp+Xba74b5YJMuZaqOCsME5/bsQoZ3TTRP
BhiJk6E9cUrH6sVSTGhVeBTqkRSTnrVtSsPG2eyhMLN1eKRP2P4yqKf7LXcaZQB4
raf7o4qdFGF5FWRnfyhYGV8vl0YTBPDBC7Ltpa/2reOfnJWniX/o0Pw1bka05pc7
qhEbXvo25ypg39Ow1b4E9RuOYqvFwGoOy0w8VEZk9Dr0eTGqVWsetpBjtvu6rg9y
vP1ZIbpyrTkJtAyO9KlFzT9IefTKggvCGXbOpcuiePPMt6kxmDggvQWfofwJXyFB
OiJmvk0uLIZyrlMrjZOt+Jh8eMrOCxuLY2xUVB7La5ggav8B4VXNlFosOGUTNoGd
8r1hVe/GNUbUfCA7wux63T8IGDDXxkOF48+SrIHTTqDAZmvrICVvzdg/Df7x1qj1
G0iq8aY2Es07jxUNqVAWrXUWtWILTbo0tdT4U4+h97rFm8o6A5PJHCg9KWPYFuNd
WQ+nM9fbwCtZ6S43qCKpwi/z1cFZS+QflOhsGXobKBYz6zkx8dNgJn3lTUPNPJ0Y
47RHsK85x4pXUT9yf9SPSrza/5JKwEzUmWcY550xTomeDBN8lDJ/KMV0kRG63UJu
x84GFCjeD8lanWXxvbriXurqwfzq6Xj0HTw76OtJi8MMoCXYT80DprKd6ck7jDc6
TVKaL1T8Fzc+DBIRv8BprF72G/5kPZCbtocMEydu5inLi9Cpxy8crLwk/318zw79
WgZiXdDEb7h016gMfYCQh7Rxao/8IBQHTQvk/mLvHdNbiiX87ycRf20iXv9x1cjN
h9JVXtfjtdB5DT7Mz3QUKDb3+RDEhJ+WoLmHaRpPr4imeFzYcVvbU5trJwTddKVJ
4qU7hQ3LlIgOoCMvElxLTDrF98AWoXhzqgFZJHFA3HUZ+UHb547YcsJDXIkUsXix
ESddkAnXMa5tIgN3K3BHyRLngX9B6CLkpqHNANsNBFt6eV557LOkOBvbVzivTklw
ijTwic6pqbQVOl90BnhfmsALN79k10bXQSGdWO3cU4SAckYR6OLCDFzdwO7JetNf
OeV/wJdAP9+LAS2zD3HqJvq7T1DlZO8BuaxUDc7zrxv8y//e3oEdU64+XVGH0fwD
WCp1SDoFYH+xlC8QW1M4cXhKfNUYAKfdV2w+iswx0K/K++sfrzfFPs2WRsA/rpI9
EYHAQsshtQvu8eQCipCZnUJe32AxY2eZUOfJ8yarQ2/SFpkXA+j1fdya9CWqirDV
PpF9VRtZhD02WGbDhGqIZ6+cwTd5+E45QUQ7Dq9Z07m2LvUJvDcqGGwSWao6RAE0
7mEIt6gog2XkXGQR3QshDhp5/Si0F4jkw4oE9SPP4ccH/ct8DcHhD0fzG1J/8feh
YT6XFXGNRzmL0qDozzzL0Exb/Ez6yt7eSDwSElkpDyIIInimmlmrd/dB8pkvu2ss
YuhGdfjmHVpsxL9RD9jhZUKlpxi8ONP4G0wFeGrpjutBrdDbRNON1ZaCElbnI2qq
M09PWQ+IidH+T9qaHVAw8FDboK8pFnUOqj9MqK4am254eQl6NvMvq3ZeOihPetX6
lKqLuUFeVnY3IBhNoiTlDg9zPZGI04s76i40ioRbmRCan5aAsLa/vtcziFgmkdmo
gbCM3rW1uwMlTAJYLM87C2kTW24BNcFVSlW7eqOPjbgPYlPch8utCjSmCgTC5JzP
ksi1SsqjZAXXw1zrOlX7AobqRIUi9Iwhp5Z6BuDXEuGxW9G/dkgokoXI5wXFfani
e081tVbMdeOZIIxxfU0BEaZiAf/+NIz5FCditn5y1wJjOiUiiQmcVc4Oa+O6V2vW
1dgCkq2Eam/8uuW95SKUC9KuiNqip4QZ1WmhRJy2QT3OSL1Ry6jH63JTX0+zLbPU
ZDbQZXtAzEzQqSizdOG43YuetsdqyslT5lXfyNti4VIdT9NuITqEDpNspBSoIkuT
R5RH+MNKggEOAhZMZZFf+oVmfa61n5LlF8tXk3NnHH+kWty/NEzrPL4xXVHddKPQ
qofAh76frmtu+ez1PD99rTQle6wcf1nXJ9VxND0NveNN18V+cGi9RGIRAeSHQApF
Y/xJoSe8hTdjcaSKbel09swkpPKRYfd3ejSs3C44WN3Nv4k3QaQzpFQ9m2ANKYhZ
m4vS6f8PCqZ83Ecn+h0/7uh9dajPabv1XSoL/q9JXNXJVV0U270Pj86yP3N+oV26
JOXlsdoc5L+8VutsuYsLBk7uathMLia07odzDQGaMQe59gkg86PdQXvvZ/71/ZGQ
QF8FD/wVE1BGInaWqlN1uePw/4WN0a0MhFW2yqweiN/4RwMXC47fPWnOxmWinaP/
nOSddRiC8XDckWeFBw0E4XgDLEANcyFgd08YwZWySYjrhhQGHyJmZQHfAIYV14+8
CMTXOXvwSZMQVGGJj9f7WCrgfvGEI8XkjQfyGbYqDhMbZuyuAXpXrD1uRbHgYO9O
U0froG38lmfWRuHW9z4k0JWdW5XwM+k+cWjQybB5BxHPn7jjUCVnzC5bzCcastw7
qeF0y/drInDKdr/0eN2ZjUeGxdm4vyx8Fkdr8KHdKusukV4DjJ4+pQBncCA2FwM8
TCGG44T9FA8usC8plWTGUEPICwbE7+kko9QUS1ISWpRpCE5zVtT9+cjK8Eto4a39
ufl2A7YAblpWdg4LfhRq5fRdXi20cFDb7ptmi2ZhbIP3cWU9OydUz4/Ab4dQ+Vsj
NkxQH0dyXWljEmd8vABtTgy6mjb2+iCQ/easEaw/DjMqwmImKllZbE5cdjfcy3cQ
c/U1eYxo/0/VMxkYE80hWfdS89L0o8orJJ1PK2S9gB5bPNrDkedjAo9ljgKyMOS+
rsCdp+hSzVqM743AC5rTM6OVyyFCi1ZDXe8JQtbWo8W/rgk7wO9H6wRBAFAmvvaO
u+I613pveEjzamWXj3bsVBBTht0hyd5+AnEPlzeYgahMcMlXSnKi4+DjqyYOxgbs
8GaVSIgGFivOWLYGTfv5WyoLaC8oncW0Bf7FwdJZmf/V0MD9cC0mzAey59uXf6eM
0tjvT81oWHBcefV8HssToevXFZBraIx1g9KZDt33oe2yfe2RqJuDnP97h3ok/5g/
RTmnT9QOqErQwV0DDLIK9OLEBUOCugPxdL/eL6cbHIfDRjr5QhK/4hQ4S+Rp81qL
Fb2bzTReBEj+474p/3JKyhiorzJn+xIbvEyRT1iW1UN/GvDbk9kYUULMNT5FJ9aB
vRhp6dIUb7zRzwtR5ZUU1lv7L6u7ThMuPOj6XBtP1G/SBIYkLqhlbYGQapGbyr4D
+J70n1766JOhbqTs70vFGcBaqFqgJDCSlz4iBDTASxNg0cbipIYPefMomaBjnp9P
4hVDpjE9hO3LEwDnny557qkYGAuuhPhCETjPH0IyEE+xLJ6LuMnCj+qKYk/5yfBA
bdsYg5VGxug7KsX0V++i5J8ZQ7qeeJIMPT9qvMGE7UfCbInwFj9luwu6/xZl58cW
6WDYY41uzPERyVfPEyZRW+3jFRVJMYO3SXPeGE7M8Ac+cg9OuZdlf94ikKPhoozd
AvVviNCqzph6hn8s5maiTeNlSQzqR5GUKT6zcAAF7dgAKsDihNDeTqvJ2reHwWrv
0vkEfB4Uq7CTyf2r+QkeAXeHZAaXmVvzhoz0aBSgqTUdDntVHiag2QVsTGROn6Hb
4jduLIEtwG7+c4/GeGcFQtVT9H91xerval73iWzJYWUzjkureCJi/G3G5fQ9e+jI
9FNLzZ6/WMmYi6mdEgEOkIYRcuhjViRXbQDID+qDd+Zge54Iqf+6cxf+Ex8tE/zX
JCkFOFV8MbUgeebiKSxfCmBn7PgAJGNwKBUkQRH2IQlmzMamjkgelDoTS5ZtgWBX
BHH6oMg0Job+/gxAQRMcyA3FUu8yJtpQ0iLaHo2qekcT0N0bn/xHUcbZovU33DCq
WK47rjacqj+IB7g4wRZcbrA47DQzuW5OD8LiV6Dk1zkn/WBibkzE87Jr+00cLUzF
ikkR+hoxRZseGCPJN+DZLp0BazN8pkHaHdrXqGBR/9bMdjzX07tE2tOjKF7YIGTz
pBxC/wdHMoOHQJUOeeSCYLTnLFdc/tyGwrKzl4pKYDOxsiCwi7Er6rn5DKyRV7Kr
Ci/3JdCKcXF03IWGci6Z16un2iv1e/BQFxmOYNCAdixKbc99AUw1xFDDGcpLqPXc
U69mNYwZuu12dh0Cmup7OplLFhi1QaE+436tfG7gyLsCMRN/69SzTkCIWh/ywt5a
b0p1HkZU79itP7wvtK/C37KGnsxNc4xMTZjvr6XnUDiNIhalNGZN/4ippto1xlCs
YrWf3dyIsvcgDROMPMbHHes2WPGha9VzwsthzED9MpbvDJjZ3DZoqq3ic9Fi/fs4
bxPcvM7OqQAAR+o47/hDFjXKOaugms1pYFPaxHMg9+ut7ocpXWZ/E44ODDG8/Zb1
exitwOvhLRA0/RcC6Zo/Fn27bMq0Mp4++tpA9e02E91znza1CEWHB4AhnA0WYVa5
CVRD2rDEM7QahibSzq2YGkgIVDo/GaVYae+1yUJ4Hf24BmijLsfoAecZTsIXQ2fN
HOevTWAqvnK5+mE9qTmG/lcrGyd+9sRZb+W548ZPGneqTq/kghlmeUef5sbz4Zub
elJhbE0Itk9nr5OT0GwQOiMKp/zi/RreltNcqNHSbVFlM50bf9nUceBjnEwinDQb
xg9lUdjJz6yYM4KRZMEaSb06xeSFgWMX0v/gTmQjaHuV5P5iiN2+1zBT3meyQNB+
0dFrWYRB5KCqAuSFpxsPqy/l+DqLf48ltuFlGT5aZNIiXzqWT8kch6JFzJr3k3ms
nIY7N3xHbCyOpnE21hWsdBxI8gtMpntFLDRGsq27xAR+bsnk+eTyTJs9hMO6zhQZ
BZdyn4RymqimSFXESGOmCRN16ByM9As8ccYRwWSOebPkAXBII1Xjup9cdso021bR
/eQIUIQtwA7Jnj1mKZSW0aODOzw3o9u7mgeHlEKujWZFaXZD5LcNa+tLPcsc+CNp
6e2zj3AeP5oIS8Uzfsw7Ll0UNWBtTxuIusKm+ZU+nig+cIXuHfpwoCW6iv5Ew00f
X4vgXhWKl8CTlMk5q9bcEuD1Gp+2RI5CTcXvYhTtTHa0kk4t/gImfJ496z3oa1i4
lFc0SR5UfXvsPd3WYSiOagILKLSe5YPLKLqDnmtZstI42DjHMZx6aXyalpyrv9Sf
EiGimo3bG1PGvd5P+mviY6ek5I1xOlISk8lBpgSaZvEtGuOn10WxYMwl3UMoB+rP
3FCJihCkRg2YvS1rU4q1j2j1S38DqeY/lCXxHYipBFgqmEM+6zR8920k6UvT+EjQ
r7vgc+E5McOjpZXws8fXNxS2hXw+Hi2ewdPa1pY8UME0i57ekq1NVAReEEjXJL+Q
WKI+hfmN/043UaFvY94n/rQ1p/1p+eLzsNzDSMEj0Ir93H947/C0JBdE+P2jvN+0
omT1xMxCTJHhn1OaxF+JqkoQJ4R2ZggVxB3B1+gTXAtgdu4TKN5bSrK4buPLteHx
h0qdAi4GGeL/lAVTwZ76lWb89i85ERtcV6SHGw23C4C5n81/M9sFDNdaNi5//C/n
QDQRxfOfqsU3ztp30v15A59Cn6C5njCbHp6t/3fjDFv8Hg4d/oBF+JsYgo6QHMuS
rLECpaHPFkZx4e2BpgEPkojAiEp7+Ub4/lviMw07OUc1fmNGsjCBzUYaXLguE4rk
8DYVOoeDpF4wRDwajuaaaRv8LXngupeViNcVhtnXvLOOFYRuLAwKyfWGpoN0XG1T
O/TBg8Gx4tsJdkL1qBMFsZJwC8JjBosdventOPpQcLdlebZpvTieBNTX8zBzH/y6
hvZsW5X1NREfJz+GXagE4avpb+Jc+u5Lbz5tm44sS3ETXFWdjXyWoVH+m2kZxg8O
3Qzg12DOXcOFfXShwHVUjT4C8SVuguO9+s9RO9iU0Xhqll0VaHzwTZjFCy0YqlLy
yxeWDz9LJEbxI/UCUMK14RVpaJslV9fbvjlUXLjav9Jx8wlkaEc9jKgEwRp9sJ3J
R81UbtkgvMfY5/KpFKBwXAiEATU8Y+rZu/8fQ3R1dO5x/gL0+9jOC1wcReABRXIA
sfjC8qlD218DWwHm/2X1e6pTwha0dEyyI2sut2ZRVPCIiFGGlQIbd4JB7LzXZcqD
mQhDRELtY2Lt+KZDl/GeMYFyDghyTz+Wo3oPevauJrQ764gxjlCbdXvK4p2C0YrH
vV/3nRPZUVHfJExuIeoHpXngOidD0wUJx7B9degFI6PKIkO5xzAgN5tW81CI+0vd
hXxwv9u+vgYbBARrmHOoiBXbEzJ/9Jet/fN+Xv4MqVNu95eaTlpa3nUU5DcGPxjN
bvuVYx/6HIM1lga318SrOF+q+aXC0lTCJ/MX+PdheVoYANvTvXYRiXBF40T+fEUx
4xlG6DR/Fm16lYPBstO6ZlEtOvVuTZuM9JBkC8fFZ0Jq+ajFHAfht/7eiTOq1wDg
WceMka02LwO2LbR7C0maqblKDybfVd+0FqRxlF83EvDNqk9uut0MCVs3B/pnLdiU
a2pFiVSrVOoIXiW6M/HuFzk+SQ5MPueCAPrxVVydJ3TcUlq9RQvEMHydluqakCGy
U3ivfNE+G8EKXcHiHbrmMAe7DrPek9GZ7doMwnjc48X5AvcEqQAqwttJHBLiq1i0
9xRk/oqumeyN1OsUh0Zsu95vgJPlzetZXIxSJ3enTC5Ta6gu2HQQAoHbHqbhco0/
lPVRN9hR0WcZnisrtRf4N3BYQMzwp7IeDusdUgJOLVRWDb+SZSCEARWYQyVEpprG
SjiJYMq8WfcEVUPfL/Z62WvKj9qmoJTv9J5lq4DXUTng6cFbJmYPZFNFQMildzlO
ilmmkqWumzdjzjqV2fON7/D+jdrPfuUvC38UBZtZE8JFUokh71MWd6GC9lgUKpNs
zCc1XSWspnLXOUSDrmyYHsJdxjlwlZezi8MZdiPs/eYrAkF+oKjGPj5ggf7DPZOo
tF4jxMQIXTGJ8JGFfh6yLW/sOd/QrOGpkp9nkQW6EqrtaEjZRFLHW/gnXpG+B0cd
DxrCK9weemJoRdSMmxS4nOy6pddhcZXsdiOJ13kuZrs83Wm4p2B/SCE2oMntUVFv
zTZhgRKZne5lKyA18NyUk8o3D9t+nA4ujpKF3S4lSlpcuYABWGSdt08JW7zVHoLo
qcKZseXDYKEx0ElpQxIE4F0eoYTW3W0wVCzSR8um7cmkVcNWLO+hgIKRHfgxJALL
hpIBPeOdHyipYvxUL7IpKp+lVObmzigAd3ubI58XdZKCVcD3p359PhoT7R4z1+ed
f9x2H1XpPKt6EqRZ4tE3ZJ//Ujo/lqHCphjT4fk8NwBWZwloxK63p2GQdJqAYOVe
euiTtgTrrT0EzMAkEHPXK3T2eazVQmKeHzNo/yyWuXhvKi1AklAYj0is7EarF9zZ
jNm8ct5Zn/JVJ4lW4TI2cBXKK78B3oMhYWfm4EbJcSBQCtKATs1RwKvzrg4zqeot
xEOYO+88ssU88Pae46jB3HLTK9mO+rz685e9+vowD8TjPCewVMHxOjcOrRtCaq1b
Em0bj6HNEcM7WHD0mGJG4HkhsROSC1B52acagoGPSymFFXJP5h2l8PPKxrmHer13
7Qu76IJjzJ1JFsplhbX0nMF6URlXrgJaOs6l3kLWB38sEq9ybOIrcsIzlTaAxqcr
0A82dti9pxN/0i4PJ5eoT0GYMNmWjgvUFeWR/nWX9kQGq9icKqM7dEIVoAp64TAM
Oxe5sNEmBlnlShwCYN/ofCyewzpeFLvpc7M2kVWuzCHsOwCPAkdvmCWCZSPc2wvS
ms3blI4YTSqDe80WSTAf+XX8ps78L0tXXyJu6c739l8oFaZ+4RdYnDmoejlvPVn1
ti0IFr5o4PIFxQxN5RB6yucnkvmRepO56/97AETHvM2o4CZBgis47i6oCD+o4VPl
cutR6WAdcp9eLaig3DOiaGHgP9AmFVFq+W7bmXsJnVDn3bPOBYHVHVDiryEi+zHS
ySonsAWFED+IN6YJ9dpPk5FrMo5DO8jRVCTxorS6U6GGqolYsC70PNjwWOsZzvzL
gjtHoXWWvWnRXZLRvaIGoJXFQ8Js/FkRkyJTKxYqhQN9Rszx8TSuI5JYI+rQcIYj
oTeF6XHOFPXtnuewDcK2E5DHQxpkcXuzdSaosWV95Wo3Cc/G7Qbg99ARt7/ei3uK
ykxkQFONQf8F6SxJNUhmaeliKBfYMDHZxZ+8BOf2jHZLIvfk+AKzNtxjwuj2EFUr
My4sM6giRuoWY3SD3rrbwyrS1wADqUBJOPt/Mcq/r9NR/xYvLmMsaMUA9I2kAJZl
Fjb5VFjyuITAbzspkGtfbvbjy6xxhwP+jd4KptTqUV+0ZOqMMZduEa/5puU+GA2h
kRQV5mv1TSsmCvulSrCnyNnRhDOFPHd19EXHmjPpYTE46AwG+ZCoLAQG7whj7WVm
L9sgNf7EL/1zlgkFO2BNjhJ+vpKMx3p5Z4ktHfqO64eJ7MwfuV3BVks34MWg0j5k
CV1pw8bEpBBjKI61HAQ1jI1sUGzJjwpN8oR+hZ3CtKJfz3tIuQ5BDFvSlxJZsIU8
YN0HogUqbVOZGK0WshCQZRhhsM0h9dBTrhWmdcnxGsY7+DAUxHnT8bsP3P6cUEBR
+Vf6kaujm/zkjmd/8tjcwyq3XzuXGzxWguTSz8d0XYAJ21EKQmCl9QwXubPRez4K
wfTWtuOfqk1ViRAenb2tNgqbv29hXt8QcaCAUVpmbMF/v2kust2RHgduDtu2m4mO
UA+filywProUtvtAqHiTQeeba3YhnXjkjXKpzeCQCR0ArH5u/+klYc08DGCsZwCB
BmV/2eYeT0NWmIoL3EMgGQ7lm9C6H/e6LDMu6eYnPoWcZImYhhxnYps4Ch2mqel0
aiYvOv8BHGgE+IZlA6M+IWTsJnYJL3AR14AbA9woCxyi0dy2ApggCQZujFYRvTeG
tV09VLUJIQnm4ogpCMCID9Ma8kLDwVxzMwQdOHV1RIDMZsu7ixpLiy6FkQiXsLj2
Y7QyZAH4LBjkqxXwBiwujKZp+TzVU+0PJqZTfJkLoRt6rureQBM0bqKuqxthnkdk
8GwgOlTPULG+g9r8WzFvEQlwxEkhFOsH2h2SJk5xW92ZMCQY21kjGve6Lo+AdSL4
u3vgXaBvXsrySMRbde+GTG9Zd8sSsLzbHb7k/2IQW4Kq30EPDlhjB4IAuGgcjr1z
HM96vmcdgfGb4Q1wqWHnhbT4Egd3zjTeGs7vcYNnyupHY5nTUIocSbcLiZQh3Aii
0Q1jXh/8LrOaYCd4U5WlrKCZ3M3Z66PtwlPA4/uRjVD3aUz9FUL6cF0pcU0zVKnn
R4VYqMPuW5BAqR+Pa5fUbjYWCKIat4b5ovlcslrG84/+HB2IBGi3cuboxbU8806i
XANL4QBPahN+aAX/k1YyDp07MPcPterzbpDKUINwV33ftnihfAr/CtVG8L4/5L5T
mG6qZKqD7EcJrbFYErxswbOJrWSdGHyiqXya4tZ0U2OGGxfq07I/sJ9ruqHTyzxf
tXjBSFlo/I0mJpZ845nZjBEHB9m779P5VLXIwAiMUJk11bteJKhdczb2lkLh9b6j
2Jzr98TYkouwBtTqCG5BIaJjFbCRbmezIUzVW420PNvpDZdsjjv7jt44UiX+oQZA
4BuwrMUSSUTv8nNcoJ7p6r/BZv3ygDe27N9b9w99JVPG8mNl5g5kaDq3W1lRX9n0
moppEi284MYH6Tk2zMd6LtL7KI7I4zIy+1HhpTywOMGIaS7YCGohCKdJMhrXx/+j
73qp5FP68cVLoZLBNQEnqjUpAAhsHktOh/kTD6JRPcr6FVApDnIEWrT7JcYN/Pc4
nI8Xg0vp64E3vyBuLKisRSv0jjcDvPdklbGL3e7fD+0kmukc+Vr1k1wzsr02GdCx
zngAA1kzNTfZcl7xXS7VfMy+tnIpTXdYiqgSBSn1Nr2Fq79OIt8ZGMQY89H7e1vH
+MCwCbL25LHXnlkExWyY65NixLRq2vG+6XMU0jALlTodN2OtGt/imVSXGogtOehI
wjqVQ7j6cedVS3wETVMXJVCt40TyXFNVBn0JRjIZ8kkc+C2kslgBBRcYrgTagFL7
X6JzWZDLTYmTsxDMuLpSaEPmAoDttO1zpr4t5yu2ZmccNxWIJWkunxrI4REcLryQ
N6mlIXbYqmAix41WP4VW+DlDc8cPhuXS3N+Rg+xmqsItpJrKCyPM97R2/ZeDgu/o
MmzQPhLyptBq+jWkgtyOz73F27esxFzzKkY6ewzuYi4KXIru/VL/MWr8WUF+K5X5
cPllrzYKzqQ1XtkxOsTTz3RzI9mlVBiAKQz3h2UmygaWOFDYjuOFEjtUchmRq3HD
mpVBgd184BNeoQydjmlOBo9r1yR9Sf9Jh3Y1RbfPNUqtjAehiiMun/Hm5Zs+q2Vy
RKY8+3Os0JlafmJHuhKaHTaOQvueFGXRVqWpREhMOOk8mrMsQTjirwyP8Ru5s1/j
AxgXfQt2FQdIFGhMMuLqqsH78O+36plVrJiaCcD0hZ3SPm2OiyT00EKR7MH/CXsd
crfzAvBKu37E1JgWIp3ddQGGA8nBpSd5thKaCkgD3o6+DwuLAlS25v7mCCzbT/MR
t+ZGS34YFbnBegeZyAa4HL4l+D7HBjSzAaHtyb3dd2aGNqnd5hl+iJi+8vYSYyxs
ARt83iq+edX7sM6MCrGkYuCsYEOWuNYDcGNQv3y86uNNEb4ZF/BDbBnwp7z+08Nz
E9qHYqAFeU8frqYzHcQFyYsqbedq89RZPJq7lqSWnxZ9pK3/KcRza+Bis5QSIqYV
+pmbavd39XLGsjFkLLG7O8X3mRwIi6PHp4rD27kVxxRhfJaZ7HBi7SYjK5XYUSKu
wtiY/4Tw2CjAXkB0WA7nXcYhsT5xXl/PKHrVU9Is7AG8qNrOP4QDL5XFO3FoPhxq
HlI8SGTsUXzOcNMHG46Ds3Qlpo/SW/VErEnU4Hva7MLkm5j1N7F3o82bSVw3k/Nw
2fgQjuchmREwNPyRlpbzkKXnjHQ3kODjhX9WAidHvgTQ28JiuVuY5vCstOtD0ZAt
kpy2GTfPnsjRCtqipV7C7CrOrrGh01Nr3n/hewCC8Ek/w6rhA6yQSY5jZKtHuBjw
jr3y2UOApoojYwOv/aVCsHL8I2PtVFXKUk6Y2yBTxw0eKDvYn0XbSd24o/vPvcsm
/ocON0nu0M4Xz/0heTuUjKLpqgWr1p7KQ7G6h2efyokXJMoZjgk95c7cjLoeni/8
4GHWXEmAlI5kHFwTNxKi1pFFYFU9my0xKbnljgTFbN1D+gKnOGc3q/G8U2pKnrK8
SZYQIAsXuWqU7MBudZ3uMGfSptgV1C0bHUkZvyQ2a7hZPizr4LOpUqnvgVMxXo/p
iDdGNLUbIopQGmKX+knsn0BRE1YLXTs99YEXI8iPBpak3YobcPkUpTR/hQ6MYpm9
wDBuje+k/Vv9YrrV9QgKSFgfOzZq4TLK4Pig0BzICXf0W6ZSOzrP/gbDeeVaIrFL
mLdWmcnq5Kk0zrjYW2GAAqjTtV50V35mflwqGSMuNCUMesvZwcB9NuUjllK93W4a
eA6VooRiEK8eQgAfJ4ySsOsRny9kEXSyAUr+YVy+PKEyihUf18ZXJ2aj2bLlFSuE
m/4mCCemuqM5nybruzwAcTQ0uaaKsuPGSHTCu3QPDUYDIgM3OUb1FoIuMv4xaIkM
1UfUusRmuGOKQA+FkTlZ6MdW1z2te71dEc5AIIghBYo1Xn0RWaMtdHyL/Gr8fSxb
AcmTl1/inYsn52sf4ccksKh+AW+gTkZt+vTSwGY1MCvreWl/A0y1VpvUtGm4yLia
LWEnREUcuYXZVLzuUCxielnT7Ky4Mot2oU2Yab5woAsivkpM8g5CROlRxA1dgcjt
5tsW5dBAUFVMZHXjxebgygnovOIOc0uptKwDLD9jGtAN3uS5xr4KphbrxGVj2MbE
m/VdnVpNR3FLhq+GAdtxUecyTxukOcofyA+SBwWccN5Zoj/x+7eu9oqYq6uDvPfI
GNJm8XOtqtVolhqUovMINgHNJg/82UUltwlVrxok2BQIP+an/s5P4nN+/TVDuBdX
vPnvCc4iirpA+gRTD1KXw2A8lZPcPOBadu2Xrup9Z1xZYvBNMJ3+30mHc9OwVIZl
aBaXVJMDw2qDnvGjni+YeYNOvZ8CbD5dXSsAAMoQOS6dihQIdWfv8NnNxdtK/JwE
+DjiwOBAeufxFSN/BR077nVxkOAgtevi/2aF2d1qN17kug5D0BC20b1+o30HIt/H
ayq+TxOLt7X9V3R1Bkkqe+qb/GcJJUYHBTqI1AQamns0OfGkIJACeAZXnlfaOrxx
VxGu8cbS6Be3CKCXAnMivmcHPpH/xUn92zCEB6KzBbEwbs4eWAcOmreN9h8ZJXfP
eArw1ShhjBBmtcH5OZdp1BlUkebwrZnqQLpk9lWjnYfKUDrHCtzVMEr2gDZnd3ky
DI9I9BD2uQIGZ892VbVuUK8B3OHFuj0Kw1HIeyKZZcmI2B2NLBdqfzwy5Whc3sfO
sZx56h+fdgB1jSnYmygsJQHjw7bZTHZprBNZrO8wHByOoKnJycx7wr6aYqZb3A8x
vVdsm6RKuzHgJgBb7E8+Ve5jlpXis14telshL/9B+2IVWDxBW7JOACQuo+Z4fbz7
RVLIwnJRV4hwg5rnn7Dv17wBGUVQprD95CIwaD+8xyI/nMH28Ur+OLA5g3sP3Y1/
RlS+sd/fWB5kouXwqrjrQ8GWKt1jirTSPpNMmtkMOnB0XJ2BzlPMqqgxrAxWKv+f
EQH9zY8N+s/pOG+ag8FZaoqFAfTsLbUoZOvZ6u3+IFjBboZDoMY9UxU5E/F4rHDy
p8kz6Dbad8DHn5vBZjGk7Hz+3GK/30zV2z6INkKpOqdNAeEGwDYMJlMWkge+t87H
Bm7/uX70MF+LyupWoS9NDX9WxLG9825vDoEgQYjZ3JbwbSNbgVKZolapr8vNP1ff
QHwIjGecSCCqAK8e5fyJm9YXooIFBf30kbcmGBS9NoAZHe+2uO0KOmK9WODJjbOa
0ysBZ1/w285+hLhRnAY/V/OIrCvdF+U7FttXdXW7IildCi5fnbfUnCEPdOemS4X1
UrsyPrNIUR9cwvCDb9Gj++LN8u0jMGr0ZcFQs5eRZJYB2Y/3BojzAhQZZlIl1EH7
Wm3HompDJtkCPaT5o6w/IzV7n9MLinQyjFsSKKRz/yL5trBnOHZhb6U4Cajl6OfZ
pcBxYCUFI2WRR22DzJfWmaLInWAz6hb2vw4lKBhw3IeCd+20QhX3Ce5TUbnveJfg
S5cOwwfCc6PYAVY/f1xu7J+mvEsSTm880BTT4BzRyBvnJXrMAq17yj478h5sfb33
BD0KQJ+ZU9LiBobCi92pudHTGKF+Qj5423MsVPKczefjhT+Ax26s4bMg4vQyQwid
vnFN6Aacay7f6X5ZRwbdw9KHK3ULNEhgadjBHfZEzeeG+i26/LrWaouc9hsZ7xUq
zB8rt6RwU9b2F550CyHMxVMYcPGHA1WzJswKqJToahugzfIMS0g2cy3RcE5FANxx
dgruFuKBk0ARqKjchVW6XojX//gtRdss2OdsRdzJK+UKJj7tVfajE792+P9xm6Ui
p3ZGudtRTXho54hvyFlCOWgY5YumykNODbRKoAxzP8NpgT1EI8RItMH8PU01N3FB
412CJAJnVM6JYCBUCxmz9YJuzp3wXPU5Nl2vVB1RSMy/Dlsw8t7AwiwqRUsr6074
p/gIxMCasZ5PuLWhqXN0XGS+XoHwOH2sm+NemAC1NfjKsWpCd4SCivWNUR9J67Mo
c5qb/z0LVCUGCfsef+Fps8AfmWxXop0hdciGyhnO+uG2vV2xl3cgsJbVKORjKiMg
mF6GHPQKSkEihWYscc8qPFCrBp7dUjlt77jppGbQLDcEVLIsyjQ63j6wEj3fDKg5
jLipDR/ALpJJL6gqXcbkrWZam1W9pyTrYCzANDWRVlu/p7AD2/xHva2Ry1zB9nAp
G4mPD6OQKfSwbL+zR9uWkCrT5jW9mUV3AheI1z61snGh8RGK7BFDATBck1B00cs/
4V/f13dCPe36Y7CKjg+SIpnsSkWzqzsC3ArnReyTkaGUTZBNIi82O4uFo/fI3fKh
w1WcRyejJMOKQBRVibDD7W1vJSih4jG8dB6i6lo4HCnjdaUpX0VOg4ietCC6Gvvp
Sjbn/nygKMqPG8V+sU4Nsj7I4+qbN7Fr0Htm7ezhzQ10S1X0dGK1hT6C8AYvxfF0
llqf1OJe+vMSaK783zU8LZ/4+WXLtRndtpmxGy/nkdAzgIvAOzoGfczKaCwLsOO5
pOKgY0gl5NWF3e1Vi+oFPRmWirR2sCu2AJEdW6GS1E4SAiofTOTs5YQGPWlffYuE
kLmm3FMYRAWedAmqXh0aE7Ynxf4LTsczPFE84dM7AfaT4ee0NpiPkKmvMXGe18jB
14Io6lxZzlZ30fABkq4xP17KYDLsJTSp5SCO+7ME6MTNPC2hnj5/ebJdOA1jStOi
Vm5YVfTdaDCSKXkbpTTbn/VDZ8fr75vNT5RmlGzqakrELSX89gIZfxyPQZDknxvF
eSkEu3H28Ulg7zahbJvZWQmp5rQAV5fmSSUtQvdvToIngH1QXHMwz7MRa1zImPVx
f4eaeA8UpS4RM4B5djK3kEs6ROvdTSECEPszQ2N6giQLJjeiB0q+uMWWZwGgpqmt
BTubKbuq6RscLtry8gTKpcIeG5+aTXyype4qFKtWnpCLESkKwpF3XewnSIkY8bI9
yjQ28YDQ6QKH47qMY/8Hh0NPWoeJlBitI2vJ8yMGx5F4RBRqAtwF0cXnqcdRE0TY
6VuXU6xj5pS6mLA7OacOn8dXDDxk5sLHLXzPvDgkP6BKa/ipIJeJ/ZgsAKJfHx6/
zVAc3p1bGpKQd4UhEUExFjuAXB5Yac+fxJtXntu0X0mI6eiyZV1yswVOyQ4Fwloe
aSrBUBAOgSs+b/JPK5dYZ57GlMVuDZbe58w8FvnsAH7uwpr37gPmfpa7Gta/xxEd
QYdHkvFlKd26r+KejL/K3Fz/xjHZxkOb8C/6QLQfy5lFZCq5SvvqmQ9Rh84MBTpM
garTb7d/XaDgfPL1GfVbd9IWsrNVwbnvfT3OR2HJsqu+2GagDTp0dfPQ2wyFEYwt
eAPVIHVYOujPTYtuoqzyMtoSleWByxEuMN/AkjQFAkC+pzssVFLcxhUrgmkrAklJ
P32NJe7WUgLqN0sJbMP/XNgRXxTkjiSGlwPJr+FyM7W23V7nS1HvfLsrnaWlefLd
NKXX7RWO4rBPjXgf6RgWRgFpMCoBBpN1t6Oz4h7OM+N7Cq8/1p1PtId1WOoZeHJY
PyksBo5d3Kirl4Vk1tDDUrJbwiYog88Ci7gtgAU1GRYPnkGdKlnctrIS53j5RkAs
dZL+tKul1RzDAGWwL73Ho30OPV+M6/oqpkbzm4lNKUM7vP/nq+Vp9kLJ8GR3HiTo
tV5HAgAIZlkDVThHg/A8bLvfcXmG6vgub+tg3lpVmXj8HTO7HpEP5Z+QqWfAS3W8
yRJAeqWopEjKm+k0VY8lSgFqmgWsCNc7DHVYxZqwjvvw+TLo/7IWhTYbIg2XLEg9
`pragma protect end_protected
