// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:40:55 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
P7i9vSAmu281I9hAAtqiPyKS2hDwwKY99YH67SGudTqtBbKRVa8VUH8FECo62uhJ
GQEvs+XOpcb2K0v7wpEx48JgrdCv4rWh8CWgR8d1eQl/SmhqS1R9JQKwavnWnczC
3jXXDHPv3ZMb6XChXAQGf3/XRiH1TGIXc+gUnf2uJmg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7296)
wuQld02CiW02i6kN0VK9eiQNUsZwF+DwkYbAMjmubzFaNWnLuYYkGJYYp/MFu07H
YzSvB+i0GHxqqnzN0wbSBSROtuy+SrkW6Aiov0RMWa911G+xwpossmOIhYZBqqMC
ulUzlqTUE2Rz8GVVZV15qmtgPWoSysNqaiagF1hYI5V21a3hxmiW6bIa5vFDXBG+
GaBNDg873IgADHkh3Dt/h0xtLAvoyu0oPMl8IJW3GCEaIy2Y0RNIRWyCb46Tk6RG
Dg1yRGEldOq0BBJP0pIdNzs7lv12ZBgpSc2kqklX/7Vz5DgT7A3vKyFHBqRPFOoh
D05ZLH9xK/+QYKli/9biSz3LMjMzLtEZod3vgeguXIdb0a5tm/lKX91GMr6zbka0
P8p3DHGkVqX2EMQKGXRDoHZS6Tq7TOPB/QZ4OIhjT4dI24Z/ogOIqFHjg0Iz7klj
+ummtLRhZgnZUN+LVrtfXgCNK1iknRZ0uZKcCiyjXp9zRYRZA5UYlXSYB/Jb5nDE
uyzW6sEykMWuvbw+103WGcj/i0GFQCfZcwG7KPIkifEhqX5oafoAjQdpgjnqiHw+
89fkHrQBe/9tfbQhoTbu3gQFoKmb4j+jOP1pz2KYVtd3jd6M/KzQprqprDYZ1xR0
JStasWiheWLKdfkY7a72itlHgytObLfszZSVJuxzc4OtadO9WfXyqAT0zK8aI5SV
1fiHlaRkhR2g/w0nvpYrsB3M/t6m89hW4dQ22DjOOeeaWpzW0CIcNCZCzTMM1+k6
bdfv75+l303Nt9annqBuQdblONZqEhFi8Zwy9tZGRHaNGLNBmaBLnPXjVkBZRs/x
oVEUnwRv62bIzSSBDK7ExUx/V92dJVskKIhzPw+T0XGqz4xeObHvHi2mcbYzK3LK
AgZ4SSSOebF+Afsy7bzq0Ow1GTPfaGl+Fh4hWj2d6wopUU7WJG92GW8VeohqWu6d
DjcTkuCMdEqeDWPweAaZmyIQRfDrBGSTWfrNeeU7V8A86ZS2OtKhrhVHD3DbSXIN
7H+1y9fWsxjDfP0hA41tI+N2awFZR6uSwSYOYJ0EZ6a40CAUVqnjA0Y0z43AkWh1
0dOlMrb2gf9voXXN6Y2zqAlbZWru6czM+zO3/DFea5HAc/+N7wBkss65nZCjzVVR
qmIPeQfYWXJVFdKmfzVeLNCu1+MVwBkQkOBvlQ0trwdWpiNVpRb/fvKsjKfQvFnO
dWw+Imju2E9MSlsN1bFYa/hcZr4cxTzEXQ5rqfzfvRDts0/DEjHF7V8ac+OxixqO
umEFHOKWPTfmeRdrjRoXepPSGyFQG4jWzSeGuDSDbT3eiInbkCXH4gQvM4yse8nz
yZqYaNZORlF+v5OFmLoHDzsnogib5Wa5sXU9T/EGNxwtxL3U6Nu/FCgCZ6DlVQxk
tHXzUljZgHVOma/hohoq97MWRR5jZcQ+NorfljuCGbWf+Z6JmXamzTGqNmYE/+YK
PPDKHMzllf8+dfFYW52vx1yMen7AnquK7HJvsBTz8rHEL2rJ7gbxXth7KJWq1Ef4
dfX8Mtl5QVD75stJCWAtGASn5H56a/YKHM4qUJJEwONxDP8p8MnaE/l9aiEAyGAv
2x2z8eRefqJ0iLlGS9UV5Gb00Mcnf0pATVO9nn3G+ZanLFQhEQ1fIUE9SoRcKxUC
TgQzlCfFCRRc2FRFaZC3JPS+SlFHDSmt4oVJoABZ+0pPTcZIqzbN0/vHLdooJ1ez
U4rujcT0R14raIsXrYl1kpAGmpbqKWFoPCEJIIGXKNBq1VgyV/f35/XA/Np3oupr
t275nitAjxxD1nDe2NVL+61j45qYsG0GGRME9OwY7dFy4uvAr3OO6vur/8mKd9A+
Lj01ULLBUtfVTYaIeEzyzUWH0/olR0S3YWeoOPpnov1Fbqf40B6s7YI5mo7pgym3
6Nzr+5GFRQj2tiQhObiul24B8otv99k0CS5UebREDTPtQKCrwXuU3hVE9nysQg9E
t6+zXt33sp+r6tkJCgEasVqJvuQAR+gME+25Z7C74x4jC6Pqgknb0NVsJasNPzEU
vwHySS86YWvmzB5JyjDpIc6AZ6Lqyfez9FA0eCIfPRzi28iEeTtd9IGBr8WCoRud
d/ngXWjNR1g/lA6l1ZXwY/MSrx+0q5OABT8v8MmFGP36NC8QB+j3zBsh2OeKH43h
s7jccfc4607KrrdQ2B5AkeYbsvGFjQCx/WLqnVwphSwVNQ0/IW6fjo5DV227Ty9O
SjdKAnBKC231zea/nfOZe0aue+Rfqp3OjwP1vRAO1ynGnwKPwIuWC1wHjnA1MSP8
FXuXmMAAzNb9fgGSHPZ1PRkmfE9HMOwim+EWyVDhNfEkQb7yR2YB2sGv+nvWbxtr
McUFikz8ne+lKooK3YelAzoWEUjapye/oMYZwVd5x+sy4AFQzeC0jJxsHo+ZAR8g
uN+oRX17wD23KQn2jTrM67dlGXqk027VJqnfHGUr3FUIpPR0AQ6Dv9IJw3K1uYzF
wBRCH2/jbL7BtoHCURFtyeceQ7oaQDuqD0D/HKXro41+Q8lNCUM7dKgIaJ0isYKa
CffFZY5oXjyEMg6gmKf3rtjWNehemIdgSuxjf73VlgbuW1R9HH2FI2r84msA1WHB
uAo7JbLHbdSMso8gb5wfDVnyFgRxIHgqPOJqosRkT/4zq94RWm16DnYN++JIH7h8
hm0PhH3pRAUfIX8PGHNUefbv4TyZQtLHsplmA8E6dA3rjPMp8BRYTNrGGTTXoQc/
+VqR8PnN4TqHgSu+eA2uN6hnTt+G+XzCLMMGFz4E89wcZJL3+xPaU7lAHTS2jl+4
bapc240XFwn8sxVtTx1aCoxWwhObeGHVC8sw6NmWwihhSQll+4FZPJm4XlLtvJNI
6QuCDk0mlphh7gxo25HVAqrtpENHgmcx9/UEXAumUPTLZyg9lnSu6232ZLzZnodB
dqMMimsVTlYLu25NBSSDrdLcgfKU6T7Nvoh1eT9YcZ1CoAUdMLNiymrDyrPnXG90
7s9wG2KY1L51p26xOuw+Hojmk/KRXldUgDgMSriTZz4/Kbxlv50AZlXWEnOYHCEm
oGrO7nBer/yuGu9FPDpY6rcNPGUBfwQRPEETHsfQkUTK4XgbCSPBY7k3ibaCZwGS
GvKn5Bm2n2Y1tKVoUiS4lFCzF/gzfh3eLztS+67dXspJCFryGEqW2o/vORHeCdkY
iU5k92GxVbX6E8ZvHN0kiKRvoTIJKk5A5elEQEEz7rfeRTc3/al3XSWyWZP2KeLk
owm8B/5fLaQR02e2kTHdxrxMXhgmdgcbbabP3aFitQq3YnazhoRvwkTbzkFW8rqS
Zwh7eIwmM167WT3kR7pxloMUnmKndwl78nE6bknX7kxb3ocy6CjkyTJ79PlpzqdQ
q/DBLreNLyMql4vjlGZwuCJAf+jZurNjfd7MFrohtF22v5IFQotpRZMf1ElZOfXa
00llbcMOD7Btd64Nbs3SJ41KfEB30p/M61ryaDoocCHe6dI/4sFdOHccs7w4l7Nu
Jv65UFNgkLhK/LRFjkbm5ByfLrP19zj1GQ4/X41MR7WEkoa4VHpP6b7AxfYUpPPX
ErxSnFFBw7L4GFKLG72VfFWX1ZY/RlXCXFKsd+Zop/7c6UnEVpxfMfqx9ooQsNqR
KFLWcIgdF6SlysxBhLxb5i11eISQYQnN/gs1fTf6yKVYhELTZL7MTQu/Khc+/lnw
fLaXQ/VhX7TO/AuP2tTHoRKodlMIJq5PktG0AM7KvkHsLW20obH1BmRiQssE84Mi
kA/mbwRpg4mkgXV8O7q9pJZWuSFH0szPOD9MC1JvLCC2FpThBCH/9W12aFN76rDQ
JUhjcnj84xV9DZAXw2/mrWtlVmE69kyOWjiueCTJvB6L5YmbKIEuqE0BndR2348J
o4AUujg8io51eZyTCs9F2J5jRsMVA7WU1z45MsXYTz3yHdwhWbJCqtdezORqrdI5
UDb7exN8k0T4y4hJ717y3hyOsa2dpjIddp4yUgoDBdIf0m9eEXfy0Bbcg4oXMaHN
aTVR0CtQeUv4oaaLTpfwOSYW/pDtGvnhvqcQI89CbfGLO0Q0DpehXLQUo3wyldjY
32g2nhVyJnWRGnOcfDwoc31hzndv5aqfv83/TiJaXdRGDZuoylEk0lYUWMqr6uxe
Uh+kpNJ/KS3AqdRuRE7PuX/8fSTtLPSZYOVI2f3i8ng1W1ybKkGHl8IpVhaVlA29
O3GCai5bl5Jayq7DfBH5BVol041Azr3GVgIbEKaOWxvz/ytHg3e4mP8Es63K5VK5
4cXfwrMT2QyL9D7D6j94y1AvNHWskfbCNVeATOCc6hmJXGwN6ylpzRAPye59Ryc+
GduzbQKYeLRpkBv5U21vjI4sWiy0dOekvbkPtfknSQiKdQNkYOhS9DDzwrc2tUAJ
Hki/OQJwpUVeGen2c8JHnSAh9+yfCkDRUAlqICL7iupSN+QjaibFm5mxKohd11SV
wymZIhldbd1iVbVjIMXbvi6zEZJo6JJdMSL5qpOhcMu3P/kXqa9ifIhAQr/v9TBD
kaEfJVLANCfyAKcF2x3ZVpzGey0cFIljVQTKJRRDRZA992vJBfnCQU8o4dm15jGL
5ma2SJS0x6/AoFBSmUlYM/qRz5iP4iQs2HruIPCY12NtYNScMhrpi5A8VHVeMtng
smBScehFnJChPkdgeQcRj3rLB5DPWjeBFDORXBorGI7H8ZUWWRzXRLr0wwzdspkQ
IBJo8wRrL9shRbk9vAGrfZIGRsVyAeyNeRIC8FXjjWHxFgzfS4Z4EuxHiOZi0t8r
GpozyeSg+KQxXuMM1g5Klv8zKl6623N/5NxGYCjDfkk78s9Q/vT1FAO9/ppdL1l8
OA6NKg/MM6s2rDQ6RzI3zZ7gQ0A3OiLdcOoja4MsQ4mWQe5DsfnAcNXTKKck5x0O
yMHee+gTNGDJw2UQhsieKk1M8B7LTokkhyNhdQ8jrKEXrhj1kzIMmCsppfZJb9xG
F5h9m7Cgi5V6Qo37FMNGlyps4FvqrTS1RJPitym+/ykMxreOF49zTbcc5cii0psh
37GYHGqHFycS15S0lfPCf5jhKJRIl0iz8r+9sEKimegTmwjCDQfN+lkl/Mr32KQ/
YDtt/bAeQBUvX4jijfUnrf2dV3Oa/Y9KCcY1KnVJOBzWCASooPHgYeYZq9WIw6HK
cicj01zd0ll1e2E6jsPMlCiu98AbmW5Jju0cjWYXDdxdxEzTKzP6UxugeVhuzM6J
ydXsxN9ksgaUt94oG9t4+Gbk34DRzA/hMYC6l+KT/9+JjNNpEybtvrJCgSmKL67t
8Dn84AgJ5JHviaUDpGnZvgE3kuMLjjYURZJdoWOe/XY+Ij61zUL+t2XiewWRvVn9
00/gXUaTLSupxlLpewrQbgVOz5LpYNKGVPpr8DMX+qluI1XYeLJ10jngcpVVGMAI
xyFgm/eXU9rbuyPjuMUELRvGMdaxHH7RT6rHOKUMxuK4auLgHWsDdCMYIppe6Jy2
jVlDAjU7xuafKIPtfsE1UeJdekJXPkoXDuGEDlnPPD964P5DbLUntS6LetbBZ+Jv
ogLVXNJk5Z5H0uPI4qKDp2L/UxyL5dU2lysHXi4sLqkRq5Zpd25QOwbr8FbGbFaR
E/g3rnKbD6ybrX15C/pE9EScJ8GB/UGEtsouyBdWPUrcHFLJu6+8F1op9Jv+mFrR
nB6emJZp1XeIzdFfho9RFBu3dOptXpuBwFM01Krq/0ecSngHUibVQELxNHevRPAJ
ODSMGQpJakcYsoI0vTvPnKcf/tpdcO+WkWaOCofH6zU630cUxDqiqObquAjw/bkH
XTe5NPgufHEIMkgKrbb0UT1dz28RBu+IjYy0kAOKxGh5hw6+1BOYPCTjvGCNzMrE
N/tInQ1QCjuQSvDmQq/vp+YzY4r4qw24FV8gknCZV6ebnD0iwHopUafUbrAgMS3a
305r9sTZ/Udb74uvC5HIatXKZ1Wr1gcbk4r2Z+UbpBW+aK4ENCK1cNJzvwk9L6R6
lVuKjzC0o8QOpWyX68BnQTxUoJJLRknIlUZ6eOOJ0IGhZ5xSJU5nsvqna6XP7jGl
BSj2pKLQEPUl2QFEs1anFjbPL2xbsRERnc53cy+MGo5QNs5v/jRX474jQoo1EUDc
MhQ3Nlh3jBrWVFkA1Pm+VqUhk1cA/ZqIVvqYS2npBS/DtSZ0xdHstsST42PS9Rmj
J421dErGDwAgBqnTn418JhVvtpR80wHuW4Zhmnp7ZTCh58zj6qOfP4tAmFWzlsky
XL5LxEUyxIz3uH2aKUkUhJPhYg8KZNCkTQ5JhPdpaYvOxzQ8aX6kfDJggEiRZN+r
S8wy005DNgjmkwIpbS9TNsA7mZ37rYYAjyK0REd9wsR0vorAy67XpK6sdtWYarYt
A7jsEiNuFPYwEFoXDVeGuiZdko7234KsW6E1OA6SSL4melY8AJoMluaEAJxEr4f1
hgh8VvGq61wdACU3/pMMCvp1EmvFzLn7sEOpqAK/zL92FxyTsclVbQXGfnYb52J0
aKxk1Kw9l7h7k1JZ2lG3vxPZkJEQLlxHzyAkXfiDnUbULoIhiB0gXvkldwQtlG9Y
pJCvEAC1oX6U8EV5xcD/UHK0Ot/mI2dPtp+RaLYKzwVnErGIpV8Q1dRB6oDDWEMy
2bY0wQe/zKgE4w46c8hFXI6fjR+JWZwPO9wcj8rxS3Sp+NWzaXAB7YL8yszvW0ys
LoWsvU9bS993X6sk7cU7Qd6t2AlepkjrdyQMgyxU82P+Ec62AumpYYKFHVl20/iP
UYdsQtMWrBuit7RaHUsFOTd43sU35etZyPr/+xKH+mdZ2SQCYTD4wVOX1lrLFGAH
0e7Lo5WOqFHzuIJa6/+xOWDTJlGNYj4F3uzHZzdGH+hLJ4vxeZqxXdIgC7YVLEgz
WktDXd44x2qBPf2OW8PGZ6R+BCaVsaCvQ3I1J9hEJmnmWksNKDPG+WTZjgIWsRVy
xfnrH4r5VLaW/kANx3dzeIatt81CxTPBTNBSXmWxQCFVduMqKlLjlgdxf4vud3jA
ltz8i8jdMl2D+lof96xO3jiPW+LVH50CAMDaCa6rJ+DUH5XKi5fuimIsDOKRYwot
LS5d7X2SJ661WjZ7lGwBST38Ygk7+Q6ZmR64+GkovTE2SdKRJ8wdcCl0n+pTOR5x
/U7+U0TqgoCPN7oU4OvHN+WXSdpXNxbc4Z0a/MG8ab1uleByJQuMqanLCRMOnPvq
UhVrrz1ucgAkTQnUFYlgtBWtv/dWcslV6iMt4R9AiAep9AEfmZIVo2pEVv5/0Q9q
RKVYA6BYXHlOdJtlK82J91R93ogSXaUmT0vwtc9zaKU6vYmCHGwjigelsPqoXgyP
a7jnuAKWgr/TxPF/ZYs7WJcY8k5SkamwnxH2iXKjMNCzWaFgq6UnyQwMFEcKX4K2
mWH/V5F5V439JYmx3O0cZ+Z4sExhQ39GxVVV4SkHrrrhdKz58IV4mKMbeRiVzDmi
ugwLDogDSSs4E3ur+/xPR81nWaJ7tlwxWj7v8c2ujDuzxjkUkH0hRy1ko4zWx2cZ
s/dNA23hBe8w4zi+vebisN/bSp1JMBEhrDcXdTBQFof8eZRFon553pwiI1F7MoS7
LkToLEiTT42zzmLEWn25ZEvluGK+ccMayeJc3iQOxXvaCg99heXvgeLJ+EAK9COd
HiMCKvWdrVGlhixY+v1stfurYYQ7m8jo82VaincTtZri/zmCrgS01yuI+LiBedMU
fMpD9ZfB3uniUfqkZymatnRquDEblqrvENXo4KVN5ORkeDFei4ODipC1XqEytD+8
nnevesPaJVOzqamLclI+hrDUgaB95oadBHzw+l7DMkJSysFyIa+vgbeZy6SnZ/1T
7Fa66Wh27Yp4tHrYvIzhx05o4PlV4DLEN6EcHj8tVl7+jTrrKzymAwRr4McHrLJ4
sSOCNYQGSgadYLACBFiux5SWdh+x+YKx/sgG3PVK976qPw1SCdBdzZilTHy34Cuf
BXNc9I3GR1nAZ5Mekwzh44TFWfY9Lv6aQKfC65tvfV/erRRIeFurkQmGMEMmN/IT
aasB6NJN9JqdtMTXRjBWY//7m3YzhG6EXAYaj8xE+iWV/3Rxr8uHex5mk9TRV5RG
hMJztfYcCxMgV2Fb2sXUxMCRcUjWradGv/Cx8WyEQ2rnf1FCmZ/v+JdoRTc2JNzf
B/eikq88n13uEzMFu75hL5RYIgxQxF/7bPNSI0vK9USggOvj3ziR32RoBP3AuGQP
bLuT7YdTuPWMn+Wb8uYmAX3hkMNZKa0n6u0edN1D2fqI5MnIxS/+x21nUbxBeoZM
yXjxhwm84zl4+Qv4Nhd2ZxTb/dDtl9wWVK9U7x88/Fr6r6QgCg9tL106mUczr1fV
wDvgaQvutnXKaja3ie9BDaVKbyiMdbhX+kCnstm32jz58BBg/d5h9nA3kVgF9Zvt
tNGBGSNyfDUYYKdZpb85vNnX3BFWo7OqN5JK6GvLD0zj8bzdHmSL+gA+MRaXTGng
GXCy+VBVXZUglYD3bNljoDCfBLZXvR/lJ1S0hqaHccOVnp8B1Cm1W0GdbSD6qHlo
HyV//1UnYyZU8QTStwiUqi2fe3YtorjyZbh26zFghkyck6qm+oJcNopH2xTd36Hz
plIrJQNaW4sgMcmeOx5MZ03XNnrmichdAYgAh7wGGgFkxIwMdKJox9DuCMA24y3n
M+9qmN6PB44IKByHhY9vuootb96qZ+I0jS68VUj1sXGXDMWV09WvoCGsLsqIF2uO
lwohMKefnSPAWE/zmZkg7ghF44N9+48yMlsw8/T6T2tbF4q9mA1JosR9S/p0nmG2
4MWA6X1lA9ufrUkLV1laKUDYzRZUTOOEQvZe7GWQnCKCptlv+sNLKLHcYcui3rSZ
bA2wDrzBIAQVqJ4UzU43sFDmmkRGOgf8gMC4SuYsUYo3DjHaOp/qLOKvoQPXX7aT
KaguG6UKrUEfB/gBt6j1t/Fjmkyr4gzM2SzWaZ8Kiqf9Kt66T7Ni+yTv64ZjAkTh
Kl0ctbWhwaVGzz4oaRgwDwniWD97ozRg6/K6D4amrpP5sjAVbIcrRUtbPhLCWH5m
VIiuTa7mQC8eiS8GQQQAlUoRHvk67jv1vbZANfWP/YpFXtaOvUWl67gOxyu3n4ad
UZ+SEqns9OviBWakml1eyN92o5OU5a90WDcA3gGEIpk1MMSt/URZzit+zDUis1kj
H0SBEKatu6t1YbJ6utd3ekHFu4e22hJ8221Iy42dvct+25GxpJ2CUe86C159cCC+
bmEBqz5s7M8JdhzgkDcKDnKbG0yWI0iu+hxOElY1FG5ZONiccoZrg6jYC8xltSFx
a+YMm6hzcBcj1IaaDSZaA/zbc2nAbj2OWJloczZzDv8KJG3PQYLQNau0Mgeqk33D
ChEbAzWxtmEcO59jTl4qBwzaA+yiCVbXcI0Mv+9Y9Ls6F2iMXCbUw0SRf3I2Enit
r20vJUz03AQ62GMIx6TxyQhhjd96dvfXOl5j7fPtTZELshPcOmysnp8bIF5iAR7r
vadZ5X0OWW4ksqQtmMpzMGoXBoqOfSngv7WARuDVzO0MnsqD71lOJoQXbMl8c76D
EwNC/CZCXTd8E8O+2p+PpWh5jTVwEFsiqa2OehwH1Y8cyWcmMg4aAfagyDVyX0lx
WRrByvolCiGW2/BTPN9QYOf2OMsvWkmX4/np1F0875CQ3LIAURCV4Rmx1ZA7/E1I
`pragma protect end_protected
