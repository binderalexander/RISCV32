-------------------------------------------------------------------------------
-- Title      : RISC-V 32-Bit FSMD Core Testbed
-- Project    : RISC-V 32-Bit Core
-------------------------------------------------------------------------------
-- File       : TbdCore-e.vhd
-- Author	  : Binder Alexander
-- Date		  : 16.11.2019
-- Revisions  : V1, 16.11.2019 -ba
-------------------------------------------------------------------------------
-- Description:
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.RISCV.all;

entity TbdCore is
end entity TbdCore;