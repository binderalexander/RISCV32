// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:40:51 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Vv/ZRsL+Jp8+DY0G39ihiMQAHBf6qRTyl7B5en7CTsd760aEgw9Awl6P0M9cly28
Sxnr3sVv2Hg7u6plIISLdo7aTuEXCg5ezh+jCrmQCyf5SAcwWly+366CLrSPb0XC
FUK6Rrtfq3RmZiwLNC5GeBcD3birGCrFJ63/rElc4us=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20304)
qkwbGZX/vmcGkxp1zdz/6UGXD/N//9lGlU/H2041D6Ti0D/Z8AyzepbCU4wlJW74
WRDxhNWZfWNGtA//xS1xsniL/kuRQ9nCTqQjl5HOCucV9i/zynGiGFOfj2Mz9flY
YmLmYHOvGqK6rxGn5Hn+zE3ccxZTxV69MYnISNozpQmNI4FGjeuz5STdL2qSvQDT
RlqHf7D+8ShLZmwBWIH0dOHwmVrrJCKxRWlfxYFRh7UaplrzagzLWF8bi18LzzuZ
Hb5FarYSy8k6amKUp7fDlhF1ud2UVrtr+F3+g+nv36ZEtbSiOEw9tqyV94ACFag5
zYTTlcgx0oJkfyurCP6hGEEvGoWCGvZDU+I1orWJEmFh8iQ88vOUZkxQ7j9fPMSK
Cuf7kt7RWVEvD6f9Y9PDOVcIXfj/N3cRt2CQ3PiUBs+GQIPxbfnIUhg0HgrT9xoV
xzQOlHBQCyNEDhXFfTNLy0VvBeROrjykTPJY7T1zAsbXjfw8Eo/xeGvKqW+ClNqc
pn3inrs4RGGAXJLowqwPCYPMJ5jxdnd9oqo/RDpDjAsAxdNGeHzq1fE9/CjgoSBK
7J99+U0rl3pwOUkSfu+LfjYG/gBSgU+39+o+CS0ibN1HBQ8lkvQ7qVKOQJxeOFpO
/Z3e4TeUlRKOILG1Sszs5Gqorcd59MdLG69Jv5iK9rzDyalTaI8+QHtdJoYoSRzQ
oUafCYzW/kwFdpQ25UyLfIUy82BiAKH/2tvOi3s3PVA6eW8+tym2ruPQxkAlwjWz
3+asUsdC/jY/Ur4fZGrYRgQengh7Xj39eQyz+dCUXBx9Be1MgUIz3Chp9jOvsRPw
+LCD85KmzBMZLwVxuESCjFCr8giu1+LPfE+MfZ2LUMVbUskj97TSFMFI5ctAS2rB
9AMn2sODmpYgSFIWgHQi5vmcAsejpMgOqSacopTKc8y/gQuU+IOit6h58ycHbs3p
8VV/ax6o6+z73WjbIQqt0SP75f2vI6g8/PPihDVZ3MkZZa/BhzaHIB5BV86sa+Hl
jsqMBSwbH3t1Z9ULgCYcNZzAlXK69A4vTfpH3Dhy3+Jl0l2muFGgCmkx4q/2UQF/
xpTNS5ndoR0dGzXBZfqvGqvxznZPsR/axnAdDRcN2ZjrNsTBe7ICAMu2TjtVW3CJ
2HcoK1PV9dSNZITF6MHCuG/+9gUNc6PQuOcTp96n/HudFeOUjfb1jtCbf/n56744
2tFtY4dQOOFcXIdqJ5OY4fPKec7p8jS8Mv0V+4R8jwBP+Wr6Ea915Rj8wdvxP5fa
zcGoWqtR6K/jw+BL6/tweAH7HPV76AHtScOmI/N2FCsMsda6fRwtN38wp9SF7AxG
xbqQn7KjrIvvbxrzenxDMoG1snz3xyEEeEfHZq5mmg443Hz53HQvT1N93jF1Mmc8
p1h407h0OjlE2HwGvmqlUOmouhN7L4jU8XOB91Lz/9yTKcn2UcXQf221IydzkN4v
wBmDQkFh4SOW7RcjCKIM0U7xeUYAWpZrxSCChTw7lqZGP5Rre0Ve8QkHFk8NcFSC
rlbfZSWVZplnY8Owmuak3iyhDGBduTVawkOXZ0f+p8uQci1MQOKeOJwbuVwlIHXH
puB2VZ6O9UAaGQHcLfIdmpUuJhc2Qydi73e35GCHYStTJ37beLvyccekHLLEpg0l
Pj6lM3agvK4lyHc4+/2sF4QTgWD2cVRejgyTWjPO+SkPLNgdNicf3QORoeRCpsap
BRDL7mdYEolNEtQ8tppLBDo4+MQACNtgP1qfZwuzY1EIXUKyjuet9GVt6d31KriW
H1rJN5xRr+7xYg/pTcNjEEW7RX3TvefJPxit48x/9l6TDeikrl1Ty3eVMb3ab4No
O9fwUEIutQC6sDzJNSbJxkMHAij8lr+ffWyyz6Way6Vy4zg1RwN99dYutmxQpSk9
wEwE02xXygg1HBSrw9lLY4qtvFFnpHa2zWe5RPrWtsUqbYZqwvG9/dtGZSXIOko0
a0o7POeLvKvWv20wqKCHGClFbCJkwwqbeQ5Pt7Myi1QcwVqLv39A+i1+tdeBuUpq
Ve5DiWfDKzG1XEtckdwWe15J0s27XR9rHXrESKFbqCIZ86kDacmOQHlsLYJ5Bvfg
SdBpmCSn66uj0ZA46lXuxS32KhUk9D0JmbR4MpQvcV407RAUVkPTGc9VJdpz/gB5
P2kV/fnDpvmiqoQWBdPS8sdtW8nhCL8M8kQ9ug0trIC2OJtDPPOrni1gib7e1too
y0yiVOXnuNha0ssBKRgLzIHkLZv3JruHgSM3VY83UPLuYzicpaBi+3RMihWI/5cC
3t6d4irVDsx8lHONqbNIw2I2TCS6W2Pre6IxP1juC6jzdJgGOscKqdRNKJR8OQ8J
18UKVUDk4O1MVkzLFa6NU8s0rJxwqd/+5JblQTrJQvk14vqleuVc5P1FrCKWZFTG
/GLoPXU3a1B7bv6hCBRvArsq8XGC+nGtgRWkj7g65cSI97pDMcrVObtGxqQKiIYq
Pi0v6utqdcccQJiVk3sKdfwuCyLxDXcvyiFKzYqvJu8oYRRvdLNa8+0zwlIzrHQS
NTcKlawMTFTPk6oZzw+iMPSj703485b7IkO7UDNG1QEGWuzagSEfTV0FSTtvsAu5
LDMz3pSV83qCFRfgFw8VRq+dasdVs4cvmXP425IlcQkJmIGmZC47Zqv+kLBsNFz5
+BhgAOuij3gMD8fxPAaNs7aLkNGdDx1xGper9h6FwhEM6ULRwsB8NKjNgKBncUCX
jHxEBjLnv8jH6+VZy6kFT3ktcKREk8IG/CQOm+NaBoG4bkrxDKK9G+Io/lv4QLNa
xz5mQCs8HjjJ18fKhSrzzbM7F2V1cgO5Pfn5lP/Ki2wS9kfJdlhQfVuqjMSSEeGS
02tNaNPXKiRVBt2X9UurTqeeAU02Iy6GGk96O7IvkB+tEz9CdaEreCkDrM4FyA+V
6wj2GX1gZ/z2gUGAJe9bPZOy/zciisRLiwK97Cei8p9jKHOs3uPEp2ysGSJJVXd8
4CojiC8NecT6vQJKAwzLU0IZib0oti4gUIvH7G8cFvhKRb7dfN3B6OH4FK0jTB7n
RSLNLFoMVNrGsGKStAEGc1tTSRXU2GAjz9C+Rk2l42P8wcoJUUaAHk0W2Zd/sBEi
O3sx/DZhjQGZAXoKjMJhrRrXHr2qndSbuYN2/iqEOa7HI0UBvPC7bu88h46na2xs
Z95Rt/30YfTGZInjqfTvNSzxxPw8gCqVoPVKU6f6lfV/5O9iNVHKUhNoylF6AbyR
sj8TBFL6JfkTFwQisEIxmdTgkg7j7zzhBAcTwt8L2/85juuUaR93nFk50QfDsyS6
aF3UEyxImrDkrjwVk8nWLfIRO8OJC4j5wtgV66PXVTtQ8Mddnfjb7+gml9wyrPjb
zQtabNsaitIACifEc9iKn0vpEtBnm5Bs16PCobsYKfznbz6IAZS4tGHEF1e2P5UJ
W9fYD0QF7O5ZsvWvZ4O/mS4BRwrtXRE6ZztX5uolBG/49oWsNwAlNNNgoGf0A/n6
ft2Xu9Ek6W7W/gCO8TFG5b68Z9qRBFSd1gzO6I3YTGYtI8MnGcA8A/qgKwTEdEPi
nuxRxN2gLiUgRdtK3F3SL5S/JUWMnK1N8bv3kGGXwCXELr0eenECwBPsSzVBsqqB
d04FPHe9LiMpcLTOJVkKeD6OBuavctUi8RLGkNTKZCXz6/x8zDaq5aEMRPjHnEA/
jBB2RR5n8QFkGDr9IMpXsH/v+9q7g0GHY+9e8mIl1PXiMVnGLYmbUnFwmK9uJSGZ
DG+HlcFV0n1FOeVAdtGurjBPlk1qLkyAr9cYiWdewoHDnAu8I2X1R+5X4jEl07gI
SF3ifxkaI1zSvLkBtlpfVbbi+2aG7iRq25DV++kOrkf6ViMCiNil9xoUB7wy7dPo
5m3MfRBZ1osd82LLJJ6tFW00EVF2WDxCAHSn/vHQwOiYKwf4vdYAYEvH2Om9Mmva
ZQqJAAp51ZjRiAcpffuHO9o2G0bABmeJQWk1uNeoi6y2CwN/frKzT67EkzJq0iKu
f79bCpK5TPm/yJOTWFXiUWIAMshKb3t+kkcRE8LEkXBF72Q6gkdOtwe5XzqPJba0
4KJTxhL9ZArRSPt0QLNKZQLrGuHUQRLmj5ZQrzvASd5DSg4G+Sla9kpOWGyKy+a3
i495ZNKIp0dLw77Ui/js/+YuYron+1Qc8KSQv+AbkKs9Koh6QRM+psKql2vvGkMI
ckGHmUTjAWagCxJkqEvL2UMgoI7xnxuEDKqwGx1pet+oRIgpGERPltPv7RKr1Ofv
dtgGoGaw9g0+P7v5V3Qui0i4HV/+SAZEwnwytSNm8QEx1G011J9trQXLMez4FSjM
q6U5xrwZ4HUbxzKfIJ+pN5TLuT0QzZZta1Zg2Pz7U1VOJWygrVZHgIDQDAl0WNnD
9koUZCdVpBn5yRG1VD/FwV1zLSGGzyhz5682i1yb/fRlWqEdVM6zpj4txgl23jAN
hzn6IliUCXrU7hWBWOcMvXSwsFuB1rhnae7yOSYZ7diN662HRY5VptwV5s2itCxM
fASBqctf6q+AwwyXAy6U6ftKs25rogoCOhAQ/lvARtCWdrhRahBlSlePqcR7uCYj
nMJVIVRfOdyHoRcaAZJhdARzn9BkhhqVnRvrEbzlflxT7KIhvnrB9Dxtk1/IR5SS
CAWPKvfV8+/J2iOAEcHFrC9gQ554W797e65zlzCT8CH8CvVBFbofZV7vZjTF9rfK
V4fjrLhiC9hvjxNE7Mp5C2vww/CRDQSfdmIGfqPw62EEfYJznpVgYCac97wg1HHK
wFrbEqDd/3w/vIYwgYFt6ao36oJCCZWEvMdQCo2xRtwwz99Z9g90zm6ao8pK04uZ
LuBM0vWLvebiNEa9J/iMY/mHtlhTh8NcuUaBzvHUimylUCkG7VogcUHAEe5vbUXs
NUSI5WGegZVF2luPRUnZrb5+x9V+wcCbBHEHP64CmmTq8w1INEwCMZsrc+eZe4Tk
xXDE0ID7yzFUEfzrJcALXVpTvH5GhMmFiTmy/ZlmMhpKAEkbaKtRG/q5mmPM0g7D
aF+feuwVwMMWwNTWvx9CQ90RDxrUuXLgV0T842nQTcjpFLQNPriTjjWJ8O8luY4O
gsFKjkv9YRY1kNsz/MSW1+4Xspdhk76OS8nqj61Ne+/bXeUOWTUWe4CZoBrLUqHt
nm0056bKUuEAXQKV2Ne4VGSlafbtKhDprn/nuLslbZTupMNi1pOMsUpu+xTgA5jG
iZMxHm0qVfrC1uQD2Tl14AeSaL5yUbtNfNGF09jm3aSwlX02h/gJr5dekVMIiNPt
wcqASrUvL9OTr6s/93/yJjpM34Yg0wuUPpb/SEeSMnDIKTkmPTJ7HSlen6gH9ylw
YWhNdUUPT/FHHTrk2feCy0ketzne4May0VivYdazxB/28KTRS5ypEZs+WJZ+fP0k
KEo/mmOUBv+JUJiT9o5eucH1TCvTxLfuWOFbxX+Dmtze66ixhFH5nHhG0o1bBEM9
dQSei42LV2BSmLc9R1xa4DH8KG1brDV0AnWJNr5oPGaqCib+zZbbPDMIUP6/bmvI
reCWCTtI+FOKWhgc6grve6Hz0eQr+X1fWR6BGavvw2+lRd9nbMqXGc4jAu6vtsIE
Ydjc7FUVIK4kqrTYFszheF34nXiBn1JpZpt9/sUEOyiKXrAFr3xPWm56OhfMMZwD
UlscBPBrTBne1mLAeyNIJU9b8rBconPu5pEwh86GElUjNOV9UKsH58NKoMFAeUv0
tVJpKepdz8LwTKeAvlWG2kMQRGipbgOGRj6NadUIOQaj3KTq3A4cU0udgmCjrpuz
VcNobSlOs5LuQM9VESk6hq4lSJIB/A5tvP5GDvBi3fnyynQfDMIdV4R/dcbCt++0
lq6aeW3AgQlld5UcbLvLjYM9MWz6er6AnpzkCo9A/avpIE+9u/eAMs4kTHbqV6Rr
V+2eK5/u087ozl8z4mKzqKkJqLiwvuFZX0k/hqp8DPmUtH9TKzRGG6izDdIg5p3Z
jl4yBKhcHGSPPF1aGZKgYzTgkkEU4RsQ34O8e9H/coow+8fxo64Q3VspshVQWOUJ
OVu9V8JuR7WI1TJPfhIwg3pBo9VyDkSySbMIOahtEe2QMbdhOUbUrJezpiESKd63
HcYWcJ0GJy49bO/fzzK+IqlsNOn8ylA/BQUERDOslWEHJEdYR3I1SFMqbCVbl+C9
yhxwDnGo0MMTZAghtOkez5E+Eov6ifKqF1CVwinNhDhjXiINugOEADwnAaXNcC5F
40X3cR9wb9FnF+/Gng6NwnRK5uFAqnIKf17BWS/Y3dFtaTujwcEPJrt4it38E5Ia
ghha1oJgvjdgWe+Ex4cHWToJqBFqxBf2K8sQg0REyDIk5KBkMxRdqFwJRQd/M4Iv
Ez5V6oYFLFnpbniTgoi9FTIqSM/+QpEk7DIO12jSe/RRYpxTx1a7CU2zQ0bZ5hna
e6HB3zM1UDIxmOSIkLpIe4CU0+AjdUPmcf0ZfhC0WZAEOcXRygemrFsAxIU5L7Zn
Mmm7dPbuIsq5VIAQuP7mWHRdaXZuxB6M+h2MTdZxkQJD6bjrXpBN70mBFkx2Dalu
ZTxAiype39hR5FVz8MVqyLHPDVa8iga0QCaBrjDSKOd+S9e4tDBW/otgjPWp4FZw
QVV5BB3pHIb9bOsC4S5eQzC60mi5+bRn4oaA+zMlf0mFnVsorSWMVXDYaUdMsPZj
RS1FPXBlKzka0abYi/htVT9aFtPxTHiApJyiRAcbMq2bizAV0GQW4tcKjE4qUiKF
kvFgA+kyU+L2bkkf+wHdEyNSe5IbDbmCzKUCWZPxabzHIDRJpuZlq3EWflgr3btp
tL/JW/uaZqQ1DVgGBaR3pMQgRUW9Wyb1MtNubZVbnrTvzIDv2DLa0+ZIfCqx0DfW
XJ+wWPwP+u60TJYf+XYbudwbeskqXRN08UIuuZrJ8QMv8uiDN6N/Q1tqxxAFGmF6
eFXVQuo9g8MIvmxnOMpbj4RMe6C5g+d7/GlfDT041nI2bNiovPjwM2NLMfWb+5ZF
UJM2T+ZI2uEgya3HJcnQLKi+hOUb3pJcD3bDU0JMvOHU8VZVO8mAX8IiQZhxefDZ
wau8L82XtRp/0Jy1ed9mIvkXnbu4mQm/xEGuUwHio13QAIPPlqLBEx1T2Cn0doUA
5LC1gaPs16oPk31p9UJ20FzIC+xdbUYXXrSiSw+cNBb+BAeCpemIkUCWuefveBOJ
kwMBrmjRs45UYTu2kVAAK/FIkzX8geZ0nrH7cSb++anoeegEpYMUFUz9JBoCmljz
ZpRxP7dtP6WCVhfEr6XgzaehSMjN7arMRBaCAON/GBz7g3wxU7izWZwlF+kcYI74
UVv9/8CtzEQiTeZYRAJFl/DRXg8usMDkTc+lZ2M7yJVerHC4HUuXV09IN+UHEPH7
l1lf6ZNRkK9fhRhK8QyMqaMWCUs+u++yztsaz7WM0eNDhBFzogJTRf+Nb2aqXj+V
2xSvcUg0xYK5dJxoei9TaMNmhNmpEtd7+yrRHJKd3aBGJadZTqioEwgl8fas2+AY
S667+WZ42RvIp20n30Up/xubz23xsflCJfeUUYrWSwIAeXbOl6BTvu4OJk6cArtY
zOMBRTAaO5rm+iPnBQ2UEs+xOriFw2ePQcQl5bDKA/iYDFo3o4It6ZiKQ6HMx0Bl
oI4T8+HUnQW322uB/t2Rojox3WA7bpDLLeCiNK8IAYSX5qlWXF//ZeuDttvKPZUU
DTdTt6KigolO7OZD/perplfRtX3Dz3TbSabFRVa3qh+sBpTLsqJA5xIJ1Z5QTRmP
nI8szgkbwoboMS6mwJHFMr0dpATHBcVT51JTf0d9ndLfS2v5Hppp16Uqfv1gkTl6
5H7yA6NNIwXZn/pEAhzBoOmcqykXfqRJ67OZ3HTss5rlYzT4Muo0UCJB/CTmC3m+
o0LZjdE4TKmICt+Tv2YyTQ9E2EgAVPrdnCVpmEifC1GtTdHpAZbPfKET92Zecp3M
OlllSkLPLYKagpStuJuvlelaVVf7v/lhm5qtStHGRcBiEhQm8ktV8Ku9fFt9I5Nl
T2Cypih37e/IlpPzk3VNg6aYyFftvQyFuLAbuOlAtgnZIeK9xAuaqxZUPUiKA8Fw
+wIg6ODvSAful42g/I7KONAFr94Pcwo52V+9Ek8YwKw6kjVS3Bztvgc8cMX9LDWS
KJOHGxTCEhxsGFgakBMK3MzkVyVJ/mAL7/teVEXEZc5/q2VjwKIou9Lt/PhmgvLK
JJ4puVy+TjN2vkdfcpYkdxz6Il/yCWbo8nVNIih/40K2U2PbfK5jnbVU6p+QlXm5
KKa5EiiBsRChTJ+Bc0QrQL35kXa/Jxlr3GwSgoNNo9RLcpAMf/ZHx00OtC6Exqx0
8PU6ps1/2nS7ieuzaBCvaK5Rf3suEVX/zqUKiIn+u9XMS7LEOpRZWWePfb11l2z9
73503o91i8ai4Y83mKZw1iOc2hkxd7VljssZeBVspMEGmhmwkZgqr0dNj1CzCAQF
8SJLnXprWF4nmIa6BgAd8d2+XsuLkeSsC8sJdQ79NkInSym7i3/83dIhtdBUx/H7
L9l5JhvaTccDL294XQLJ1Q6Qs2UJFFPwDMGVacDhgzSZ2o5DFoLLn04yhPC0vPjq
vzFO/jsfBtfl4kwhUMQuYu0VrE+IKIVAKlRg4eSp6Gdxz91G2HNjHzn7UAtKkrDJ
4l33b+dtd6Q44wjx6ZrHdkmeQh+I5voegE9CBfCAB2f08evjJYFO/yAW3DpChCBu
lpH+Gv1HQ+xvC8fFo5ov8XcXifsmqzjr7jeMT5xV+dIYwQbBl++SXrLmMzBGYCi6
arxRVMQo1aCNOWkIy3mmaAZ3gnm+C1b2FqpHxn7JBeIvTHi/BoicTrrhyivGZYEZ
9YVqmtxMgt2d4bCtXfZOtMyYt+tvRpM3/JXXwtdvZhXQvQJOpYQKW/JzbK4CFY4I
IaXzVLi+o7mBG6qrmTUcY3dKDEdBk2AEfN7NfeeppqlspgHWmZd+VEI99pj6Is9O
U/keUICqjFAsJZwHZbAZyUks3rYHUQcDsE31QhesH+1Aax3AMzHSGmghBFr8rlrv
oQDxxsi9Ah9B06CX9WnOVKNKtxFZLW2ucJu6+mtiS0Mx6Ru0QoEpeJqVi4yOTEWa
ZB/eS8eOjJA3uxLzjUpbxeePJrDdh8VuWsHbFxYgy75XfHM6zxaxKHrkE9ov9avd
fCiuXd1hEtj0+k0J9wYJNEffGFNPfdgNwnBNcpVnJ33t9SMBRKyvmmCZtsqm8zkC
hn7GjQGJebdkcuhmn5YUzPJAmzL6kh+y0cCD+rqUs5TdxSJrvZgx1X6Y6GRwwSGR
BchmRDp9VCT/J4l07Jp+JpynOcztRVLaYrUgpc/3TDiynplv5cvtPOdXoDOJt4NI
pt/dH+v81nS6dYEw0NhlY6N+0K1Cdq4FmEzpqde2H+eqXYP5nuGVOiRueZ8NDGno
hbxEzfEZFhvmPftNXVYDOMblmJN6tjArxTb9tdGcXkJGvZpXazoojpMlLwmhH2Tu
680LD8wnkrBoTnxlArofYa9clMyUaK+KEPzAOZT46D4R11VeYVB0z8upZxd3/UWt
XAvJyNppOF8BXXzkk839bPzOPqmsOqGQd5B2jahCZRLTAnd0mBGdro0nAUcZo4qA
1vafwQ1bCFb6wee6wKTBLpc1zJqDcoEY7a9oiC2WL6RpY9GJi3VOHm6+f2CWcRTk
v7xWZ/9Fm2KjKYLQ8k869g/DoWPVsvZucTXdkwa55/h7wKJ8BKWuwDgW3nehmnKP
qgcbgBMBHtHzP7Mvhriffw5qn8anBkYfVZQe4P5+n8wMs03ZfMt8gtEbwMtsDl4W
MxtP9jr59iDtmkqyqoP6rEh7QebFQVnic3s8chh49szX3NJRcsvBuvK6TOJN1xZk
hytnCljerqNk89s68kSAvL3EcyznNr9NtvPecBGSdZnikSDfbIdOa/Ylhi/cPW/S
Yy5L0J0t9zwHlK4FHext+Jhkv32EosOZefCspvw9BpB63AHOl8RBOIZMrT/ll4xN
cYALn7nZXBVqZWjwOFvAh/QRThPRxPgD8foy33H/04gm/PzJ231swb2sIsyyQjg+
N5QySwO5+jTvCv1anc3sMNn7V/e3PZMrMDAJ1q6eibDEK/kovSbUln4Yb+lKbNuC
FCXeOmY8Z7nTGKPG2UReaDL5VP6LpkdHOL4yKZyZ90CpwXUHge8zSoiio9OR4gpU
VrQg9iP4l2tOp+cSlReU0dgibXO13sDtgzLcL3tCK4esDol1ZAWiHfcpe1psJ723
Cdh/OunarJWzdAW3YVbDCUHtz/R16NGecDV72nk3Z47d8tpm8EFEyV1/kwGbe7+E
3ilZ87wefpA+cU0TWYS8sSzAIM6afJHjUIhBcAAGsuy4j3VHDgZEwpb1qxGIZN0r
8SCFouyqG61MI5FQFChm/K988gWhjc1SLFUZ7E6fHPVX50O9Xs2yuwvFvd7Kta3x
qX91faYSv1mMH7WS0le3ymZ7hB2XzmAiY8M6vcfqI92qhf65Hj6cz5arc9MdEdDU
OkORg0ceAfaBjQuhyDrnJwfD83uvlVGiFbpsFph8dBqnU40uE73O4HRX2TVcuEVl
EDQpSd0CQduVXTnKxBn7/U7ZSPRg5+p6TOPZfz5yhL+LYC7q9dfPauSpTqx96z8m
yHzygorDYNdWBTFibvAb0PwymQ4dEzFF2KiCvZtDLeR13EeudkQ7vvdubJmAB0Cd
opxFpgi5b88wUAmsAWUR7rinPtCcyepLIUXhMM99jNYidP/Fk/za1kIhAeOFm4MN
uMjl0i4rEP/inSZB8ysqjHw265YqozmUx4rvBX43+zUqwDq5AuXKGG/M+idPSfJI
iRlhxITX6y5FrWryKF9x6VXpwT6qCCKleI2QZDU4bbV7j0p0TAmyTVNQZv/wVtwP
g2otvMuhMu0upPLy9QMamc2Ig8j8LSLbxmH+HLmSuVYxqCTXr0eAFAuF/R4XR7z+
Z5AB7kaI9pYNAuJob/aXasN6BONha6YcwE31dOGw3fs9MFBYHNoUZXVCyIpWRXe7
iorHy093gDBkYTDEd2KIkJEDMCENZDx18shOxZYzmr3FErm92ef9DyGp+WWe7hne
i1NRF01Yv5oOLxiY5g/83UTUfseFfuWL9T2YwelBGgIcV4GW8q4Hzmx0qYp3i4o3
bVOFPTvKLhFGFFDuY76p/nGLgYtZpE+XiwBWyqvRvLMCReg2CCai4HCm2572QuKE
jVGNqObp6sySHMzmxCyzSDhGieLwcskAFzkjPjaFi8YPJQVL+fB53xQF1KfZ01vX
cMZAq8NskY33QsFLlN2jLsg4Gz/BBGTm4oJdLFS9ofbbKjlQ7bz+sgD+SXIYhCBb
Y5qSHDbNRMfTKQejM1qYiNNRGKU0hCWqoziQcBL1T2ROVyuDWFFJow5dc4+yKAXi
OHY+LAmHbX/LLv7zLQRKgI0zoSj4kKjfIJJT7Yw87PtWCumsrhqfH97agW23kYLr
Sb17ytp7w/2p1/xhjodIG4AMfrrHa1BZcmrK7pm9x65E9zEvXhd4nPK47kF+vpT5
DOM7MN3C26qXx1APXa+5SNMAJgNyrDtvmilRL2Tbfm6owwg1sEwrlDstOcCH9Azp
gVFXScG8Itx+vfhaLF1cfZ94MMf+Z9P/pIpG+xKN/qb7ehch76m8h9kIM/dEDOy0
0JKlXhaDylx+jqzjLnfTqRU+Ba5G3+et+jFxsOwwoPEYXUK0R8RoJn0iO9Bqawus
ifG5iVbxqiwFRvclIEVRCp9S6+hM335CC0Imy9Uv6eNIq4qG8iA/aH8JtxaVJQh2
4DYhKlepdVb03YPfcOK+o1kg0RAihlFPZEbWg9kKKtTUTRXFmydqAXceYui6Rkjn
JeRKRqeswhbDqLVSFcLV8WD9jKmxXxdl4fXnr3qO3IT1jrao/CCShWOHvLk3evbk
AIcNOwWjYR/4XgWynr7fPTtjzlWvoU0RR7LjXKwldIrT/mKrt/b/9pkGpXIPsnJh
5tk37IR2ZNL03vwmyBwKGvmq+PqsJ3JgdRtBtwTFb+r52QAXb52grR0lgl7rzMz8
ZgBT1TXkMfd3wGwb8LTzbIiZ6LEQD3B4XKB/YKG1Tf8yadzQlw3jz+Ui8pr5hEjV
evJKtH8j0m2qbE76R5p8mvWYWCxzsT/cI42sfK6niwBZw7HRhPbdLGmCmiTS8lIB
4lKl8+nb/Rzb3EMCM/O3SugtnhIqc1ttpQsce+uBSXWL87FUtpkLpG+GUv9DbQ2H
ccej8fWs3kG8TYE3fR7Pv6urvicY2HODgkjF2SQyBDQ9bCipFqL5nXGoIrVOdm9T
WKWlgpD5BfnrvuIonoUwxyZdBZcSIt/V9VdjR+zcvdpyXq5yxd9IdRy4i8V8gW9u
HGVxepU4e4K5XMxfp84RjHau9tA3ssV1Ulc9IjD7qqac7cp0V9gdD3g6DpxPZMQE
fDu+UVsF1D15+3cOuIGn53XF0mu1pUSP33uhnLG1l6WUOzwLAMnJSe3G2IpcWzbG
evikn3Khg/kobgWRy5rF9eIeH5wN/EbVgBx0NJFaxHCuoS/iLX/Ymvsd66xV3F/t
kvlrDhBTAEJoHWvMcPTLAwIVbEMdKL8rIRJWlQEfvj/dDsLBYEgw6kAXVa3xw2eE
MtQdkqsrSEFi29vSNYBDrRQ6i0V7/4kwifPeK80VKvyG1y9no+HE5BgFVPYbkvQp
fvlIJbs0mdb6dDn+68t+3Gg/WA+cRuyQcJvfUAzI3INEJEZSSUxZ8TkTQH9WuNjL
asWYI2uCL0NWebYTPAuAJ8Bn3fvGUFx9UYmMI31KN83KrwMhE8x1DkgX6Ld856sZ
H50ojCDUJAFcXLwBxvO6RpUjgwMJTJ4vNjz4+cIMhMNfkD5+YTLqppbFTCjVXdTW
QH53WDWKPgjN3kpYrQBcbbaou73LambYUGzwC+2TkcHY+z4AP/rfR2rwOZcw8huI
yVCIrWeQYUIiOzffcmG/MaN4d38ERqduaqdfV81EUYtyb44us9hT+gKTYknp9SG+
dUjmfL4uw4tN41SHxr9Ldtz1CES+X3qllAxDZKllYNbrk585r7oH8EBN1mM/n5zA
vxeKO0bZK+O/yNsEqiDYUuNsn7zgXaDAWG0Usswzh00nnpu6PxdCfmindBe7ysea
YKRDMXq7N9JRqEJWLYgIa91dC6Vi8b87KZItr+Wn4oX7kKwJF4uOtEGqIz3iXTnM
McnpKu3Bf1yo8WTYJrvTibRtgcjcH+5uN4mPT0hOgKlKN626y6D6GhL/M+wucvpG
dqY/FoAkW3SJ8vwHULLT8qdHeGv56Kw/r6oszERg4pXIDqrcKJBFUwsqFI9dxFye
Z2WvhAh81Cvj30fZjFsJ6iSHU9+IqXz9zl5cT9LhKcbWSblmrI/r06kVmZHmxZbg
vKgVG2xxDzOYEmjnspDNIhM3Z+3uq5clmhkMfjf/Jy5gjuKh6x8bI0qto8RobEQs
7A15gi/c8iT2o2uCUQcB/Yx3RFEbKnYG+uOeSSv9jh/LnFn7yROiy/hCK+1l2dDo
IsVB9CxHjP93Cx0vnFSXB7oazSUsssHaKky+e2cSUzATTdrXLGh2ZB5h9wcjXTzH
eF07PmzRGCcdS2a3oLduphcAnZ60w5Cp57ObtKNF3a1phsVYJFQezAqDOLv07gcu
JWzflg0Rq8i5gY+oBoVnHCqDi9LWBgfVx9Io4km1M1izdWC5z7/b4BhVsdKlsX0k
GBEzk1tTIQrGv1Qmqrwy2OAKlVRJOAasyAPgMdU0nBR8YetOxmRVd8Eo/6lqvGG8
P4U67TI1otS7hPAH1YIPxiM0GkeyEqt7SXJG6GEE3IDPJs/T7QNlAjZRDsAG9Np0
59tCclwvGppPhEbY7INkntVXZrZc8Jw1YzOUYF+zTWZGvbW6PopvCD4RGIrkZTIt
SNPySdg9loNSXKakpNWAeY5/Ulr6fhOQ6SG1VDhj0Yo7rrlXEo1Nuq+mN1QvBJDq
9RoVwv7ztCZtTJ9+nGpFNzFeIBqLT70vBDKiF554jVf8urDF6JdfjzSIQFgyRSJf
VVgQZFUkh0zPmEgTAtKReA3OE31rVgprXDyNUMc7e1Yi5RiHQ8IrWdDebUCT+4MB
kNjRILTm5Q3nyp88o2cWQEdESbiEoD9qfq6g95SOKAY0ZGOKstl+Bih2X2D+XSo4
HOh4pnrurF3gQ6ua3qfcEPgYqpOW4IrYPF8ZJHF3vNbGAnKCoIeoG9dxdM3go4y1
CiW+qQgdIjaYJ7R+krTpkqMaku43Z4qyR3asGWj6TevIEtJofUWCS5mXxmwqXXiX
xfhW+QQCdar+5RFTr4eZAosSR3NyMqYfdklUasNb1uovJnOi4XcO3yKmnXR8JZJo
BW+42aRZY7SnRdE2N2rfJo9kzOvc34ue4XdrcFm6Uz/+cpduYKAZi80rzK2tGDYA
uM2yWPGH6kqNJ5wZFx7tcfzVc1LexE0ovhMgZRf3Ev87RpiV3LYnuTtP6fiWkY9s
lz6AXFA0JtjJu1hS2jlWD7rg7Ao/1JHGGaAFl4TzzIxkquQ6v1FQii6L3VwNbFJo
DwP+2f8Cbfp2cjbNqkVdPvmKm+yQ4w7AfAovzCW5hnLVz/BlZj9HDMO7qeFwc1Ia
DP55DXpMzDvAchJb2fXgoLjV9JluOb7UYL6j9B+2Mrk7rDyJpXl6GOdbwy4ZO4P6
WrwXG5I2YV0z0TMd8GWrQeVQscyCQllyYOiuOonujvPLrpi5rpYTYRB+3vldPdPj
/4/tZOQ+OZLbaHYkDNR91CK1wFZuiBHCj9RvyxEMLXkqNcIKMw9X1lTGI0HfI9E9
MLavbQzZ/pKZgM3RwIfXSa3AS9I11LsU3gbwvycYbSokMw1mCoMU5hVVggMJnHNs
GRCFKTFGj0JmMbji0Nlp0XHajaFbrBdX1hvGH1QBeHnPqsFcP9+gi1csPu6KYWx5
aW9tyXzsY1R3JxPbeNjRlREFsrJZizoHougldVZQqIQ1Nd38PL3MNbyWhEakDujc
drjfaQwSMLEZ/C6AOqSirRxNGZhI101k3kyIenVI3fYSnxKViOb+fCOjN5LKA3Qw
H51GjSHJCo/apoWe708s1GUPlD325yp0NEogStEMWeRoyG5eb/Y1Gy3AXB7qdB5v
p/22v1/QXfSvx438/AFkpTjO3b8fkmYL0Ux1kUU2mLFbe+a3FA4Fi1Zll/12RwyB
uZw0flXJgw4DH382QxsM3GoEaRMX5IcswIDgVUdhdYlV9pGOF26g+3Tos2pGwFtp
OUc4P5l2UPPFuq+T7l6jm8q7O3ujhtcLUD2CxkhoYkmwI48q7Ehowt088qOumXuS
Dlw6dopOGshHkmokbdD6cWC1GSrnMDtiB4tb0jIKJDwXEpjaxW0odk66bHaBOQhp
f1Phfliq+Bq/ulLkG8TNWGDhKyqca7p03D2AVbBuZgLmxZ5tJK28UiEuWxeDReZk
G+p8zMNJMadeINh9Z5cq3QE21hqT7ogYjoYKWOiohCzY5bd3JOQqzeJPv/Sf5woq
lTFKEFqJo0kl/Dul18iX//F7HItZU88RZvhlcxWt1qhaNqYw/z8a/4C+5RjaBHRl
FqZQoVtkO/LfUTs3LMBaUDo2qw6wvZiqH5OUyM1ZGQovDTyYPYSTZadm9146NXUH
MfJy2mK20PH7hkDtJOSQdYS/zsP+Rs0PtkRIDqpHGd7HtSVR2bcbBDVDxrLm55s6
oKnMWv/9Cwz72DbGWDTaxYjpv5ycNGJlO9GtwQOpXxbaGz+iMs02AmN3Jq83AiyW
A4wVXIDPjEswFXoZAkBBuwjiSIkxtfRwc0RiwuYuLrJ95nkF4NVAZybW/yUPArFs
H+d6EAR4o3FD0Q0k7XBgcwB/ByWBTdpD+lqvAQ5egz7xi0G38GjDZJLBFcnr6qeP
jZvj7Q1aBWJN2MQcJTqmQMzL3odclAzZTFJuD1EokFM3MR8p/z6wjxQizT5HSqVl
A2RrbDzetRbAgxBZNuZFdta2OTojZ9LbbxqErk47X3urMnJEUKIryciugVea/T6r
eZbGb0U/KAjV+ZmaivT4LY4Q14seLD47iHiV+5bSOFv/EE8/Snd6L5vktTy3ZyZG
PQ8Hbsd9tmaLA8W8A0fgwXDiP0pGZibz9Djqv1kZZAlmOF4A15mVZqAyekr7B4YZ
HGxwx5YqFlgrQMWVKrpS0cRIExZlTdD4X5JbKdGJZjueCMqq8rMA5DGCmkv7Ep3w
/LS6AoxJAbUgr2HFtSaWWelxhWyw804OptfniZ31G65yi2xlqQQ7KzzHEWRVJ9p1
5WGIzvDQ3yYkTZprSHfMwyvCk3i/gQTHnd5LFTaNCZiHqkKs4dmvzYTcrOdxTsOo
GXlV+7TIEhpu6GuDkUQmBlKt0zBDyEdSlWFO7ZLoqwWZutVboDifEXsFIeEj98nK
j9n4ELdap2uc3fnWpRxKJxmVrW/WWGUr762oocq0SJaNgGKARhHx3YySDhgQ60UZ
Q+K+3/xh7k5243TnY5TOeG8JAX5U+jcnP2SeI8yOVsbgdbCmvGcO9FIfUqrNtR7S
MRwTRbVLpW1rQQyWX/4EXbNWI8cc674/9GvykxxD8i9Ab/3gKRDi37Lm24+MhUch
1r/PR3i6i++JvAF2K+gcEDfl4fidwrgdvduE4bTyIASa5ydb02LJnOTWhm+TI+54
tcI0qpBOli3qvH/8Ilb7wbVTdYLqKeU8vUooK+Z2u056q2SNZ0GOjZf/4Ey0jSCG
m69vDMnF5+uvnUwLRU9XO1f8+GYz1PEcxRW7K/S2lIoroM/rMeybexDgI9u00QvW
AjYpsSp+oEAru8V8cvdL83Jb4B1ugpxkYKGcBhZCSjZyXF3ubyowt7z7uy4Y0Yv0
DsNGliVuP7IfC5x2/9RojUri+jCg2v2sxBEcwtceOxDzPXZ317veoRafMeH7eBYE
HvWPOBMRLw5urEi8lDalOWdNJ+7iFpja8f8/Y76FhAz49do6xYwSYIEtZj2SCVHV
6l4NDRK8RUvDJstZwT2WnCFFZPOmgblSfwN/hk2ZrE3r/Y0FS9waSe3NlvMovkzA
u/WyeFEAB7vYHwaVfvVKnEvj61bKeJaEtG20HahuLmfMVLJULbUj3Tc19WcJVTDA
JB5XEzYmxqTLE9Q3Qw23/ugJWBJkUkT+vc19gUp7GpURKaz6rxaXDFM1EJChmoz/
vUAn+BQd4zikm4rwh6/MBnMQwsSMagtEzBXQaH5FLzZULSVUN0PdpeoFvlozR9Vv
aiUXF0qU255uJzLhET4t79hG/b902i9T19lqXZWb1KWHds6p/1hDojBoJm3+deF6
/DXl6YFd9u78b8CUgfLRk86xD5h3Wp+yrTqDj1EDa7QHD5ECziiwXIZrATrZw5gO
ME/lmpj4dwXlJnehDp8XXKvMPGOuDqfnon86NqhDmvQZmD85Jh3EoioFDk7R6OQO
DOf8jeJht5oD/ccRiTWb5oze0Iq1fqDswtHNH5kFBINMlDJrUOGT+GDZfnXJhge8
5hVCmvpheJzCaV+i0yeIVAno2GEQFziiwdrtBeG5yZhTlOAZaHwXOEwASH4FfMyE
A/6jQh09JzDlGPzORVIi5qh6pdz3wNsrWeSUaezXm0RRJiy7RuLl5eAWdQQNVK9p
ehJK23wSVkwTKLC4P7RRwoLV0rTTs7kdH/g04pgcybTy27thqN4iHwNKX9k22j77
JYGTgggJm+W2zYiRVkaDNPFbg5Yh1mxmhptuG1K+RVuAQFOoQAdwZgdIeP5p1jrV
NjJDTNL2AoQne4/wPMVwOH50P/8Djfhbt/EB8QmNGHlnnEjWLGNzQOWFvBq2MChK
ys6FOPwYP2G7HuM+eLMXKsD8jRi1n0/V0NEfIZFgwLjPGOQ/eqR/vLnroLlRx3fi
0eXSpBWoziNTksPrEDF4vHq1zUFH2YXIeARYuU4iE4LNTrcI7EPn59iHJ7HHv32P
3XnzKB8pkdAeWO1b5wnjHNSA/dAMVY1+svWy45VTTtnJIVYtQS3BQF1TwXG4iKqF
iK5RPvGTdlaaDy4nFh+PEfvTZdW+XVHq4sPTse0imZquk+ZlZ+b1ixvHK12LkhJt
GQYQjBmeVvKs6MPT4D8LXfXklZ8e3pWJjx8i5sJ2ool7JfCseKplJzPvuUYGUMdc
KAebdOSdFBaRjIfmypOZae8YxAZmonSg0uM4CEa9iTnJ6YUA8OF3tplI1E3sqGlH
qtA4sbD5HKenV0cO8vC4N6waCesXHfEg5XUEtjg1L3+3vMk6eNmLS5lXsycBrb8P
U1bsu4MnBRthtqJVyuo1MGoNciZoJ+fPTMCMG3UNYYDqgMinJgKmaRzPKrWdlhu6
DeWKdzx6H7gMA99Ep6As8AmeRjLzQfvlOykUJUOvdEMcsdKVbSV185JLV5ELnO5u
7IcR1RUEhVVafxvWlxNM6TrSnbVcaqEEAj1CfmxYcUYnHQpx6R5p08ubZbrRbAlS
ZBZaGm6Oztp2ZlnTtEHj41vzmVu6pV8LtOaK4O5e7WoVwuhtSrw1y0MB9cGfBQzS
PiEBZkPyZzpJgtnCiwkxdtbBtCjnoZuf+/9l6+U+kL7akmrxg7A3ttzuZgV9jcP2
gTfYNJ8TY6jIhvu1u5UoagRol+u75c5QaAqGTmHTIiU+CzjV3ndYXph8ChMM3ZGk
Nm22VTYkC1ul15adZTnQdPKj+7lOIOcBHQcA/f/12+ufatwJbnLrKCoVmDMHzViU
F5hjkA3WI7Q24D4xNyo5OooqIJ5DdSuNtUh1+Nwd0SqLIPVkVG3HcCcMR7qJlQNu
iOX8+ReNqKoJJb5SPOJrYGA58b6nSX7NfOxZ/TZD4AqXqNsPuYW5HvxbLhqs+coN
N7VTjI0XABDHnNO5c4VBWz5UklXkfltJZc0cNfkAGIE9j3u/piVufPL8lPWbxKel
Qo2VN3NuuTsbeFWq81t0NJBAn7J77Hb80OaT8F9qiOWsYo5/JDRagvnjBs2Xq1S2
8MqbJSRk3WViZC6hoFrwbFNcvSBi1yp+yc1MMu/XCX7xIqutEAtivaU0cvXEpHma
pTWD20BUhxkTZBpuD04wSL/ffuMlbBKoIzxXR2TXFSIrYghf8Pz1rMkBphPOir7L
SrootqTyLt9mJ3aPUkfpj8CLkFjMVnJtia35zoKBKEm1W52tABQyq894WnABb9pf
3qOFIFyvRCkSMqtw3qJKAe9Rj/XqW7qj9yo+qHS6k6EGVj/f7HLbvv1xl9H/b1Z5
v3ijAkW7rLL2j/nU+rCMMZSQY6LqUnwLaR4Vspgt6OlEn0QzLQqEuZc59ZTfaxuj
WFQBoop95tVKCGlO/km1M1yqk9CWjDB0IIwqTEcjqv2/MXBC7PyPuZ1w9I5rAvIK
9kq2bAI2Y+SNB5yH2QN6qp5CA9KPOn4y0hPjF3nlrfNJfNoj95pzotFWlO0YCa7O
AH05hAk6Osie5s/i3A5ke7iPfKO5p123EmKB3Oiyr8Z9cwN0vsWZvmWt4YkyvY+C
DFtqFg8Cqrl/SZhKxLgMQDgl+7k2Qa04mGnOfhabfgoyPw1tS0u0wwQvZtFPHMhp
ckC2X3xyX+YDFw2/wI82L0F00meI2GgdUbrza1h1Yu51K+JIfiY3qF5k9640JCUR
xq+kJwaZolP668KHwfqTnIM24jBNke9tRZ1Ho0yocOuUperFY4Dnw9HTJNzCNrTy
nSGDFZsT4NMnYBGTPLNYrn0ODw7KQOSMEiCmmA2u9NjJChVNhfqD6x6M/XLMR7rR
iWfNu/bkrSXzIEZREU0axPoPWXucUkIJjf/PT1UZ4hvX1N8iOldLBkWyoYPXuzjt
b5F47Ddj1UX6D0goQ1LZwWFZoD9gIJvSePy2VynwC1zrWXiirtLkwcrP6+5vPRI7
ZFSxX1mjO2EpL6KicM8oqkR/KGtTnTqI+LSxbcl/HR4Y7hxUn+879yXIt+CiPj6s
g6DRUG61M6eHO3z3x1PkcyuBrNP5hN3kp+NnqdWLQ3yH7Aigncjmt8VOsWa/jq4g
2xIpjzgHNpg+/TxN/blUVZJgjvd1slK+PeIo98GeF2Fv5wAFY/h0KMK/uOqjCqCZ
q+kCWNLHva8LFWszOSfueFmO97U+euJkFsymSGaXRth7sykH0iLRE3OrqsL+spR5
ykEwecdquPlPlgUpYur3ynQctkEXEAkWFhapB/tTqSKiQAdfJI4gIbSrQ/6VZFdy
mnJmENfprALkYeL71T/18mZLOqKOv1PVy63mkgzdfF92gm16/KxCL3A0zkqmQNqs
qoXFkXQHINrcS3IMvWjnSlN087BRJBTXwVJANO7Ev4F4OBxBLgfgmDirBo35hHBL
UxPVwpBr2yijHsHq29x4He8huE4npXUAEtM4YtEFwi7h6ERwdFC4edFfvENPHz9U
dmJQEPIJoDwKeVfvU2/DxERFYKiVnN4Kn+9g1o9CYFaRwmAA0k3qZQZgpmc8ATFd
CD3Z8yMrz0905tM4LrX0PCOlDEPECCAU974Jy9ydyovcJqgpemSb9BkyYr1gB8u6
nvmj48DeOBK5TYmm+L/GTXREKyOHAWhdTQrCcSKZYFnkBKMlA+i9oHQYBFqYnxYx
5JK3hCTdVOKXTZIlTABwg5udnG/e75bl6UoA1t3tfDijiDXT7apxr/8t4HPui3tv
Ehah4QR8wmN1B68CiyDy6f29RsQIjissIghwwSY1OjHo3jNINrxxoGnDGaqRFQYl
QBBv4HVRZTPORPamHm8ot5UNnSv//zFVOdeNKUPTqx+1M8EOa0UCaCY1ekDX4jxk
LKHpGkPfE29EBsetiJfa5jf41QYd8y3D3aXSjKYMic01vRMZ8gYMgsu4Nj9zgb1m
vJjY/ksUd67F46ASaEkfVf5vYtJpucBSIUK646wQzV8UeO3ErFzD/4jq+wru+1EN
V55CmLgEGdPZ5hmr9JdluIBcuDORZuyxCTXuaWxc3tBOIG8QzUh0F3EcwsYohQu5
00MxydmVIwxICplfDUJwu8wXKJ8yZadcDYUOCEK+QhXM8LatlFplxllttgvkcs9K
oGORAwRPZTQtEOFeDjfoPbf4vC5eBVd8MO2Bg4q113anm36hqHEbcYyMkLDgqbdf
NYFrQcMza9q6sByiP8aNFyc9jFu0lRG8TfPcE9/cxbm9x2hisayWzaJhf3jBjaTH
Tpf4qKasCyxoQ3D+iOzJ7Xx+Z3Z8GoOgty2GtF4hvSs2YC/L/3QgynHA0y+w/UaL
5vvHMVApylzLp565q9kim+F/giVanqgIW3G66tM8eLzKJf2JQe/z1J3erAYx5HQL
cHPQC720RjMMDFzBsVn+Ut2lC7/zbuf0QrfrTR/u9+D5MuW8TR1C3dzLKbdb8hKn
WbrD4y//2/bSwNnjgxrHUaYl/RhEiShFlOrsfaatvGYM+Hw1qTIWJSXY+24tewWk
BKGEjEQ3yl7mESGhNt2CWKIf0UhnYUGfOhfg5/qBdomfvJ1F8WaiYEh4xbWAEfs8
0qX8FKggLrDU4Skpfi28/ivcnwyjkRDCKp1zpFYOFUlLBKkQrlUO8m8GshAJT6z7
D161zTMu4nrJwi/hna1h08RvPayyZPPfqWW/Vl+5dtagKgksTrQ+IASROZS3E/K3
ETQqBWyrMXo+3xZ97ktIo4cgBOb7YPqKkKdQg0WTQAIuinjkKCtLb79qbiDF3SCT
nHBIXen3uyTTfvNuVZQmARFceNk8EWgaTteXH06w6uTDHdO7dIBr8W1nYUrRJ+Pq
ePUGG0B9gKjJwaqig8MpFQUtCUot0t3YCm0bhd200dN6o6/dhYgckuAo6Y+e4RbU
EEg65Gbt9/5Mp81BQzG7Gu/jFx/aoFEfT9gc29qLdcDk8trmgR00wKQkY8O37eja
gaVxlmsVxWNPwHmT0v+yMQivXyr3ZMeXRiBQY9UGcikyONc2KNSeFhDTUIs6Vt7R
UJ2bzqtxcQi7ZPpjy5J1lyhjMt6Gj419lTg1nBh6mSguonJVqhHh0hUWGWmfNLCu
Zs7/R90R7sJislUnIKUbHeAyxgK2eIaulHKTDG9x+73dN3tBs24FHGqdIjLtXK7+
E41oCGrf+/7zh6gCdTfHhC0pxMvBP0Etzmjo3Pq/x6lf1EDZpMuZ5IFCYn/H3xr7
XyPWUg3Z77UkDfidTX2lkNBQ5apYmNgnaBGhoIoU+o7fDaB9sIMN7LHSC6SEQF1g
GbwgmQNPFCTkbEvzEKLGMu1qNZECV8FS3of9215Kjfb0XJgVPovPwtxBZ+BfGVFk
7gWXjAiecEJm6fxX9qUdZIGCjl5OX65DVdDCbi5BpHViVa5hbpOqDJTS4ZnPhm2k
hC6wrEzC2PIOSFPqv3bcCc6YNqmCru6ISn6bn8bbxKaRwKYv40t/mFq8uxkyCzE3
zqVs1/CnQzC0rSjPYxX4ASqTJnmyup3wc92ewxekGOjwkRB3A4t0X0LrpzUVp9zb
ZMlpA/aqCH6zwS2LALbZwT9MXnBX5QU25/E9lCpuZXbe3J2G/dgM1qrmzgNc+s0y
5EtBUVU+xTvGGgPIW2RUzyqc8uJSAgkVZDbauRsVeZN4NwYPeQKflH5B4lzUEhQ4
go+tuZPRMFnb5hqogxEPI9uBvu2e7Wsry6vo5htlD+A4Mkz9kA06iVPriNo8LO4t
nZuEWTdUI0d095n73tZHHCnSFvd1keCTRNBC5B+c2/0q44yewes1w+czQLm3cAp3
A09aOE7PK8yvwGKJ+o5yi+pXtFao+DmshW7nZDuOaFx8/Mq04TjM00c5W5tnVtBi
VEuyxMzZI15tJXrOWUG7aZCFnyxbkFy+DzBdpWe0tU5y0jA1C8yCWekEuIm8nIl1
qbPmenWMgXWk0DOVUzYVYOi9WWuMYIGJoJ4FRFEVdrMffbN4eiIt+DlJCTKj0+QO
khlCkRV77mRXfGgOt4UFhYqLiNmU88LD0jEtLgB0NiU58bm+cqFBOYu0L7fXFUpg
DzVxGhyPAnH4GcnNUeFDXGQvRvdK51uluEXX0zBny1eS59i/mA/sKgc+gNJW0wxS
8CWG9KwS9ffgu5S5H6ulNDW7E3/K/xEvS11DsgyiRwYy7MuoeROIk9THqKZvG/xN
rHXslxj1LWM7SV8shLHQiuclHT+nSw8LCD06K57cxR7bIQ4tHnVZvHepCROQBX4+
nSYBmCOfBCZElnIp98i8cdILqAtaPp5XGgxomyDVXkQbOQsVL1U9W71MgAq0FU6r
absVpbrjoiwMyoyTRd6LOF+Xaair2+JnPguaAJ4iypmBiI3iLnQDn34Hu6kJ0o3D
pcowZYf62JLjyWAumhh9Lk2yhaavSzJcoI7kNa5VIeHMqBLejbuTZylonE29mctV
s5Uh/erKaKtw1iVjYchpZzvIICDr2xzvbYFUNHsLmc80q4l4T4iY7JePflBV4prd
C5/r4vzJHxXq9wJTyYb2yDAJfW8veWL+nQFq3yDUOf89gp1FVcG1Nd/o++LEhNXR
D76BQ9iphjOr+8vGwAO3FTh5Z8lNAuTvtHNrjcOkzPT3stz3waGLLzQ9SdTUpT9R
AgjC4ojve1MYvsf5EXVP8RfhYjIQ+JjXbrN90QsJCIx15GAGIqHcYJRpEFT3QvkW
3rAnFgsRHXJDVxPjykVo8Xr5pwkCtQQpG07wI90hJRqrZgQ6pJOmxDjbyNb4/yhQ
i6r416pc+b1d8KwT2Kd1dzaTxK1URnmwab8lgrh4lMQ/tqVX8A+lGJe+XIIEWKQD
Uv7ApM+NaYfIWQug6qSsm8gyDG53QU5EP68qFba6LPFNBqvH3f86EYV7Tz6iNB/V
L1TycCJe4tYKX0oCNo9J8BM97s0aAQzO2NMf8INkulVvtXaLCkHSTUcS4/ac4G/M
XiMnzRbOK/M0OMl1eSsu6o+yc4yplMZgtzzl0QRm8Uz0gXyaM1JoPzA2rVD96OPA
Tniu3CDYDeEypjhn4nbGOSmgeEGMWT1GcOzn/6zka7pI2aIx3M5q5rA+9wBaBVen
Kgd7zVwg2vd7ToXPDn5rHOWUs6m8DOblLvH1jsZE0PmGgA29u6UNfcQK3zmRkHGE
RgRL6n5Ko9dkR6cSza9ZqbhBmwSd9WcmwqnHnKFpOX4mEF0dRiytSpMQpVIXr/+X
49Sg6NPlY6F6YDoksmeZa2xiZizZ7/jChaIilRhmWGjf+u3PxZXUnSFa05hQs4Xa
ZegNHl5qgtHDeGeVXcp51oGI3BdVMvCo2P1LzFdyoPtIuQdncuyKlVKen1BGv0LF
vaLGBNbSIOyIJ/7j3YqL45ZyUSo+6sTi1SI+C52uB56ORWGvcy/MFSDm3rmm+/tH
5i1NgTTfrT8QYrfkiMF9Mb/ZyLquQxkS3Taij8rP/K4+oe4TuM4VsAkU+WrhlNW1
Wv7vCIwbC3vvQin+xwD/fcCuO3lWggUSadfG2xzn6yPJM+2s1uJdQhHvFODMYqe6
MVVCm/NJqsTeGGwNHo9NezEjoTCL0aCxAFidNOxyS4irp3vHcNDviQy4LZnWVkS3
N+iWETU2G5SX3olbxnVSMcPXSvdnp7EYW90XBkMlUpjD3chwwz2F7V7kpGqzjYCM
dXOmnZ7n7k/11SEqEMCFTLH9Q6SBgajTL4NhvjELbWXYsPzYuqfz+0QKVWwM5I3v
U2lBrwaZbcvOQLJMRn95JoOdR8xFVVBfYtf73CxxvJuuM0w/ec6na50x2048R7rj
SPQM4FlWHLuKo3Q1W3hEv11J/vnJIyn7g7L9stMCbmDI4ypFuyAoWgq7BvNm6GfP
or+NwDQBcqIqKZV8WAOeKQQ8RZmD+2WdtaVAYoPxfDRPuf5NUGs48GEYBV69RqXn
9DVFMDDJXdUFiUEhZZ1sRA3NuPyoKkk6Vxlc/MocQmVeEz+5a8v1hZgZgnMCClZ0
VamRxxTMj5nCf0mTS+kc5yTEUpteJoOXELSzPb+WXwl2upixH1VNJWQtJ4Zn/Z18
9nYLeNZiu797nd5F1p/0XwVcF6y4iDw5t911BzXZnegrIn1GdN575zaXf/Wcr0go
g9mGQLCTop7D98qn2T6l992Il5XrmTbwVH5WIg73dBzUb6UraLSDF4FYW7kxHlct
k1+wwysIjXyOH64QOjM4KKYMuwakTcGYwcpNTFStdYkqk45ZhuEfdTNAD2H9RTGS
vM3f6M6rZGz5FWptbVjUjBd6bZSMftZ8vvDs21z9oeWCM+x/4gMpEpUMSOPXsd4v
Nm11GoDzy2kNouakxEyWokOGNR2RHuPbsAqeNs509DMFInAdMa1AmYNXCguBxNIg
UbQzEKkoa0cUyGfBtZ30CdwM7C9d/E7QGigFFcuQhpSaQkbK9TzgrjRYyh+RZwIw
76GYKhhJPudj4RNqD8pvciBT+TX7/VZ0Wqo3E3MP10MQx4t4sBBe6Yf2w4ZwP0CK
N7HFTBugMqlo5tdR7fUJQi5UeQcdD5MhoBHqDq5SJpKC6op51gSV76KKCPLadbqf
HU2o+lycPJzejM0qRMMoc5j/SnMr9s9tZWzlV3x5h0Ikhg8aXL+CleC6jcEPLeeF
khObOBBBlkWgKrLvhcW+K1o+iRZXMHjKud1LN2bBfdsSSvWLaE99Ar19brZm30TI
e3cOQNKhztsA6bmq5hUoey17QzrSIWVy+0x1KWjg44xXU66sLFDGkWlGgIL7tR9S
qHq1+PKbGA0q9uBHzhklhg1nsnSFWfjikfeaQsskS7v5P9g+GbUaRxVV6yXA/YhS
vHwm4TYZwWWiRNgJYA4nOmTNEnkvquGeIZ6mSRzQSV5Ay1q5DT6ai8a8ENNoNfix
olvcGiX6nNXKruwGzpUoltP7dZt0YLlhEyDBqqANIZeZg4dc0k6j+d03+7twFX5V
Fty/V8nvK5U3rfTIR3+FTCESsn4PeoUNck1D6BiTv8s7UjzF/gKBnJjtgn7JIUyN
dK91YGjzspfQVZtAo+x/9F03ZGn/eH6IrapTA/O4fNxDTjYz/l9e3QAOfvAp/6ct
S4aGN4pso677ftuYGrjPXXdzNbFgAMhDgvHWVXDS81w64bb35KvNSkgOLX4qZp/d
q3Uzk6R/5YftBWyy4yVixWt5JPKS5kevMXIYh4RQrOMpX01wMOtyn3s/2sFfouUN
RlF1O23WcxjMQDK1jF4U8+n1CG3PQVSA1KQ5gtNu0adn6M1lxggzVjcTlprE9REl
u9DGQ+HtawBFyWMdRLseeDJpRJS1FHezKYoYhvxSKezCXSTmkqDqXtMHbsUoPUyt
1t9YCtpLuzDuwgJc7rQxR3nB/TyNFzGqNJZTIy7MJyVBQ4OgxL9eA4oGZiRx055I
L8nXeaDVDIVg3KI98RNFuNaMfoJejbzJynUkBR7cJKNiFs5HZSVzpoMeuz7DWTt3
fIW3BF1kbtJuZCVSt4TZlZvTJbZeO8KqGb4FS7PZM0xsMg/cUgD2Os9j7FO9Fxho
0UZNr8LYyyzBW5qV9OAD93+edzR09LaYdny1Ai/+4VO72S9m+dQuatPtVn+RM4wh
wcWtxlNIBJgzhPeJ46IGvVnSZ5FmT17m7O/orB1zwAUKviMuCx251e2Lit4dNNj3
HasRf3DxPWwb2Gn3eyrb3xrjDSCH2DEwnEpKhxT/oGEPe3f9VjXLjNunpDfBMkbo
/FbyVbH6Ne2oOlRxQ3hWKC5fQ7jvUu79iXTQ9tN7SAbTKPuNYFcl5Uwwha1U5sVS
DiQKEpYzpQOIoApvp5xc6cRZlQwFnn+dnAAY4CCi0ExzFs3vnVQNow+ty8TsfYvJ
pnWK1p13/rEfcm9IbMasDvFwH2gEdty0NZyrvS1YmzXn1gk+//IQx9hyKhETk3Wj
2r/n1Krb5TVngD5XYhkRzFX73N8l7y1jz5SuPLvKcOOqvS72ve2q58Ri/a4th6IR
I1P5IXz4xzLFJ/+463Gg21fXcOVepFoJDvzs0kRWzfHmgXUB/Z820smRkrZ/hkvR
nTYRHSaVrGFB9MwZQ3TLmG0PRKpsOZA72hVVQdq1u9FwOl3Qsp03/G+8+OTSXCS/
Aq7NWObebM6AatNEDenqRo46/8pmfAqu6P6nZk62+excHOr85d4nXt663HzHbcYE
`pragma protect end_protected
