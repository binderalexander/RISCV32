-------------------------------------------------------------------------------
-- Title      : RISC-V 32-Bit FSMD Core Testbed
-- Project    : RISC-V 32-Bit Core
-------------------------------------------------------------------------------
-- File       : TbdCore-Rtl-a.vhd
-- Author	  : Binder Alexander
-- Date		  : 16.11.2019
-- Revisions  : V1, 16.11.2019 -ba
-------------------------------------------------------------------------------
-- Description:
-------------------------------------------------------------------------------

architecture rtl of TbdCore is
begin
end architecture rtl;