// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:40:55 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eUvNa8Kge3S9A1rRdMwg1PRPszwapTBlyqpA2GceBePLflHLHn7XN5J3OtNxDkDT
NGAQZtIyRkb77AcmpuI15oiAScCNsf+VCyQTMO9u72NEJNjwarjXPLUOMUuuRqyr
el7ucF4athVFlZtaf+x8G7VHVD81vSIhgeeA7WKE9wM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2928)
vKjHGfYrjVlFkZltjMZMkshfL9oQKwXwIb3K9ipi+edZJGUgFXotgaSlL+BOAE4m
k0xV+rWELvB4Xqp/xOWRxU8Rspbf8NqefkTvIwGWBR0zx7wml/5Fgs3qBtGtHfbg
hoqm+ofpU2qOQSwz94IExW9iwaxlmDpbeYHLjyiErS0w4OAAx038AhBJy6wUQtS3
UjU9lqwwDoHqsq2bSguMb1XGcc9NGe4NkSz/2HU/VGc+ln3LsRLdUS7d0uB5OkwZ
tE4cUmdopIT1VafqaCt2+TlNKzf7M9hhrpkxyy8FwPkW5Dejp2OGbXCkjapB+lpy
bLCeMR4sl55L5x4PxpeQGwgUuER7Nibgmoh6oaH58Y38onD6kEkH0iIKwHUojDqx
Nwh6SforYdobYbgsKAPxSFa6/nH52udY66VIpdYVdl4c1rxG+P8xqVaSrbUr7sIz
JvcF5tn5AQrU6gkBHBq1YsXF+yI3WxFrskNHXOnYnFk6c3LoNrOXX55349yU5+pY
ggoUGVtkSIQw9q0tEa3c2pHNphk2ju6h3oAVBd7Orw8EUbWMgF9ct03ybDrr3c68
hW7vxvR04dizcUMjTGQs+zAwdLjPEwswpYoBdlFJWXmpw3HQQDWpyYQEezG6PG0e
s73p1T1l2B/C+cgiYJDjuJhxEKe+uN28HdNUTnDBNmEdhmvTJweWFEYSP4WHxbkk
tU0mrePEL0vxV0wdnQFBo8NPEOEaP0/qUBDVVgaw6Lv6+lVhBnffJgt3kim9cKA3
U6cmPKs6PXE6lyCKkHm1PDGGKXPS2AoOw/5PuO04g3D4nK7KesGVKttQ/oiGRXY4
/IXaNiJ/reNDhpf93mQDXHMgv6OWzqHakPVXA5TRFBF+jHY/4XsPJHQk/fxioONZ
kJstyqsusuJNoqeiYvUrp+QLaTo+Eheoa1pLedBQ1vjqh1j4Chk2z8sBAM+fVDhj
F3HJ18Lka8t6CLCRmwqFOQSMhriaRjkZMh4+9n3NPIK/RnxM5DxU2dFTaG5FUK0T
nsKEVPywwDXGEkHEaLWiZ3QsDj7H4uSqZ+R0ykXdL8rw4lTseVTA1Ecv2kQgJLyC
OfbQbdReB60I1E9WY/vpODU6lqsd+bI4+G4dllmzNuFv0XmwWyaZ6wrk0l3JIXSC
m95ZUaMV036RtEzmle6Z8+pVMwjKFtJRFQ1bO1hEzKcKaeQ8WRpUH2V/zjPUdSAe
ggMrj+sbibLKqq68ljjmlRL3b5FbxHnfI37cJKqi8VyhdVp75hoGmYtqhPsiBTTv
dJbNcuVapb+A08RCU6/+RREHoN6iY5EAY0d7+sZ+nuEVSpkqL1xkmIJhvQp0k035
u2gB/GeBw5r5cRy36WdSJcN7z0dcbxk9IAVEfi6md8jYKO1nuMi6/LlKQQTppdZE
BdE5ojaqNkZ/kC/p0d/R7UAcDi/MOp48PY3uXIPthgl/fNUU+4hLc0vFBhJ9yNSF
0bnqfAlOHow7P54FoeMKnBfK8pG27qEIwpc7iV9yAoFhfi1DqFecY8ShiYCPkded
mOFDFw33UjsZAKSN/QzKFAn+7SqUIi37Pji0k5dRUMwBfLK/gEO7z/kPUnFhPmUB
O8o3RBNJqTxwr7kAPowoa4T8nD+cesNOeiregK2NagmAiEPXX4DL9JymE1j7tbgG
TBlD0dKfNCz0PYwRypgoGKacrfaV19HUO9MbhdxlCMJZBPJRSEhLOKSybD/Vyn1I
eRfGTH8Uv6+JzVZ/3KYu53dxLOLhHV1qCXLA1dbWbDz/+Fl38QPmDvW7SUdiTFxc
nUKGnOKKbb96XNCzJ3Iu/F4pWfqTnBhoV8mlb0KuLKP1gqr51Itgiot5GONUwgDU
OGHUd+Ov1tR5rs/xG3eLDCd2iNkZsv7Znf8AnBLGKeZ7huIAXhAUK6UXtCNupmHx
37ECYkgFIqivjBk2gqqio4FQstu3zEGGyyoNgpudduB2Cla67nGfVcjnHs4ofsVC
uj+gxrCdDMR9GFAADkEhJj3+nU2kz0D5Kue0CKXOBdBTppce5E8n1mo+BzWV+xkp
+bTuMjrhw0FBAxzk4bCHvgURb6PcdRUGf9hyQU8N7igac161ixd05u3tMXHqdB78
kH4mqeiSkk+DH+4crEMnoLcXDHKAux+SPXurjg4h2M21KnOnBNy70aQuZyhdZ+le
rBIB8/gfUmyQO1m4p4wHBf+dzRaAXbRfbK4fGgoZiD1nIGthJ4AXGnctWgtuh4Rt
aCdm2O/CFtHC4cGnP6O389l40+Ultq6C315EN/DexUDN3vz7C715YzNChc0c3k4B
9Ko9BL67U2XZqKhEClsyJ/+hxM8q58teG3fs5NGo9FcSxhLszrv/rTJrQXWy8BRC
jjZvK1yKh5bmu7cq8sEslSY96ZSPCiDNfzNx162V1oHhOwg8t6BAln6iiecfNYha
DZrNhmlyXXp03SbyCMF5TlfwLGk0rEjVLmsJ1g/t8qz1gq4uzUKy3nQnxaH8Hxg2
sNWF2aw2yP9nHAmsMKu30/8/hQ++DXmWHMYguChwWEQ55na76b7cJwahytK9Znjy
ZmqLWeGXplmsZGRmh5W62mxlcYTfsw6Eb9XHmIKF9tUlRa/nPQf+pNYDZLxIhYqR
hzz5V36b/5sFAuHEj1vptKWhOPfzKQN5rDmdhd16jyRZFZf+0ZcpHW9Ir1QXxXz0
lAn+cNrBiyVPlPJIDpsT9HeOs7CQHsm6zdYJHKcFej3S+k/ujU0L8IiHUpt6/dcS
vJBDjCXIDuPk1GVShuSchiKYQ4qv1ZQrsVHGU/fdh+pFWhXkUaSJDY1IA2lloAEw
aXJnlibFGF+IAuZO9VSPn6P/VSgBrv0Z0buAavnXD19KAc/pwSxIkqpFbpZb5ObG
ITq8AU/oNcTFdKqgo1glrEN7ePHKdUSwqj06TOElEnBGXKXWZlOeF1ttRsYGvb+S
vFVc66IIpj+xIFI42p4tkVVZgyNzs+4xViab8ZZFsB4Y/9FtVnMolX98U3VXYtND
f0qlhnGLdpRxM3EvS0D+zc55vsBmU2wJerOPF/HyfaTtD0jGYSi04Druo3bQXVNt
RetL8hyhhbDIyKZoJoI2GbL5bO1+TJMzuEvkFOcVR6gO3cs6Y0fPz14lBfb42TF8
jyANeULgVlPrhPxK8sVy0A9QHrSKRZ0DkUsP3rKgO9j6Yh48aZYUuq1BqCG1YfZ9
M34wl91oK5PI9exxm7iuZBiVLwFeifndY+naGC4LOgNdIamPSNwzETp+xIa+pUcc
8byVvTflGi/ZFuEyA2TMTZWfE7ZSaY11jmX78fa/MuG2hpWvguUJh3xv/eywArog
dXLC/2Zp3JqtKVSSGcNAY/rIQIjmQla2HVQjcO2n3gyg7kl1AZdVLLSVA+y0iF2C
bMxVvpFNbnoINy1Hvcn3OQfqeTPK829fw6PO4UZS7QIB0qYkTRFl4+WmuuoJq+oG
8LxThbAIeyk2D9E4OIuCVTD2dTq+bzFfF4+bQ4mY4nl+KV7kSPtklh4E1OYkBazy
EdyG5tKKYkXjGdQvE0knvJW7LHefkjEhlP+bl1sDkLxHkMafKowqPVmyW6ycr9x3
Tjd8zTEtrWIvcIfwcIoJKwKY+4L0RYeomBRUyars7R5Yrhqo0ihTBinmpM+ulbXp
e60uZVdY6vy45S0T/0BjZQMwauxvqIaaq8/sXbJNeW1hcIagMvoE5ve54xTZS/2V
D7Sqn0Uk6BP4a6X20Yn0GTSt8OJY48Ep7NW1IQjHOkW26JAZz/LXW7cHCBdo5DYm
jVQdqpc9NzYASvxlHKd5NhEJLLPP/py/YH3aiXgVG7M/l/maGN59Fx6wGYro3p33
zO6RF26SJepMmhTAnrrD5PbP9OLGF/4E/4RtIoJM/YUJ7emN+1v3rtSNEmdlEOcU
`pragma protect end_protected
