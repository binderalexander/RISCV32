// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:40:55 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fteWdJvQOfChR5zTaeHYj9FDnyqN4BPaNf+yHY5f0ctk46Qq1kH+wLuFFT0w6Lme
p33TQQXAHw2qEFmU1fj47l4/rMbAuuL+9dqm0NSkd5XFN/kZ457JFFwJRwf6A1YS
DgiQU3K107HJIHMoR+ynjvcREXIgw+Q0JOdcdIW5u3U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3232)
5BCoXsk4HHF3NnI4RqS1E82sHREEkKYGTh6uh1UiCnHjMutrOKyJ1ORg4w0pRyLd
xbKhInjnKA16xukXRkYcXeA0d4n5t0iW8Eghkx3bEwhglEjZyhpC9N+iOwWgP+TM
ODid64QkVNM9pbj9drMeY8RkPg9UbJiWRRDhxRNqBRzZRYu9Y2Dmzn07u9r4PVff
g2XOk+9AYiGBi3rrRBH0MJNb3l/mVXZhC4hlcY0q5G5ngZ665AEvkHEP1Xs0oGj5
wgjcb+y2LdrTEoIO9bdmXUQV/7Fm4iyTzVkAxOqNDPjIQeoZFqR7Ta/tNVWG/iOQ
zkQTS7BmvPodJXoETGLUnT4uMC8aDyU2pYXfCtsPHGPdhQyDwAaZMA1GVaBJLbSd
UWZb+0TuUzHNysm/GAlwgU8XKy+CPe+Zl/efTO6hO7TuHXxCUKSP3tsUC2J6KX7P
u57JMBQ5yDnmTvyGoMaIejD5I1faervaLhbbMVY91ODV2MxK9ljHZ8vwhDSBFVxe
rsKO5r4cQuJmLENfvcIK01OG+01PHo4G0YRpl3W6/D9GsQG35kUZEFVNYG8TJX2H
IymoxVRH7ivVU83x8rMVDWoH2ImczpYPeVBqf1ObE6r5n+A/F5K6y9ebcm0cKM8K
59A8TPUscl1WmfF225N+37J0adXK5F95D/rZsV8lDYQTsCsNztXIOT2FY7vLv2fO
fveIJ9EEWDdjyd64dRhYvF6WBKK4n92bi7/39bLGnxeWn43+m6iXONxdfcttgBjC
w4QVvvuWam1W/bVoJDwijpprkK0zyo+WGb0GxKmSkATv0gybnPVkDbK340TD20uA
NE9B4YFt5Qt1hu5j5rf8WTpOD1IebKhokm6mwEVrGTni9V0vFUuyvTeOHuWdhnpJ
L2uH0mBXxaCvyoP5JH4Pcmyaebg0RtJr3/hencqKl1nfwO+wLU5tbeFFIOzxhJrJ
Jf/J/T4Zjbj4l18ONRmVntOw6ZzmN7SM1+PFcV7UqnDCZkACV2Aw7OLE8WZcqYn+
vfQlr5p0UgpmPks0S1xHsVvRwcXdtpHs/0rofnW58xIFyeeGOjD7K7ntm/UrA+Ad
J/KpY/FcQSmn7+7WP6pNuAmJdwxcBLN5mVN41BwqQovlqhPMpSjgNMv/Ng3M5p/c
ssq60xWONM5AogL07dKg8tVqhWnKXsmw+hqFE5iU8updQfVUFoCUSYZGIIUylhZx
dpEr+cD1dFNvkVBtnwzJYlnXigAnEyJ65Kf3Y5+G/ti0FQWN/Qe7l41hxlEWn319
W2QK4CE9azXuBsmBbs48VuVQ7xWb5mrQV3OkCO9K7ln1AuaKo5n9F6mQbz1VWzBJ
RaPPd7BiDMgX+3uqxyGeVvcBBB1P36n7nC8PhvYQh6LEWYMAQhbP4yo9Bv1MVCRr
glbDQW8R/YU3E2+TorDNLNq90yv9t97MZtQiepbGwp5HhbiYgvsYxM1Jk8/SQtEZ
G3J99F34l1li/X7GqaHI5lb58ETJT4HqkCGBeRJ20sEBY/FNKi8d+LV2BLm3AeSv
C+8ep0MadkUhwSNHUdGrzmzO8UPe1G7aXah/7EJ0sYmgC4Dcjucrgb5oq7be1Lqk
8R/e1OcOgxKYs+bEX31d5Q8YEhhOs5Pn1UWpAa2thslEp2oCF05R3R108vNgr0yS
dU8jK+Y/VptoLSNnFPFGgui1PADg5wivlzhGMjHPCiiBhSyNB7nn9O9Rg/+Fq11b
xx6WxQLfkr8pSeJ1Rp3eI4LCYwjkuj5LCwlo1CfWTF+OtVHdbeVzh12ZsYzCwoKF
gbDBhJ/Zv1nHQGbKPGiV39sb4027La4ui4Cm7n5MFXSji1TSbwZ+BlDZ/mujRKaD
eMNdBLokrguIzgkP3KY8qrCcbMY7ASEYa4gY+nXKF4zfdaHC37sLfWBJoR1akvwL
mioPdvnBFYnLhtupRM8zgtPQjpiDz2jcbSxpvQdAnJI2I1jXaxkJiLFCCumLZpQ9
eP6dZfIDs/9xaHWOEhfeZ/GeU7d3fcRpZE3Ry7m/4MGioVnZq2Q9MLfPJXB4Jk+0
VbHg1O9SCF6UZ5IIiqdXPqSj7EkHiWJg91BQ1zSW/gSH7kn9UAg18zDKb3qnGD3M
clNN0vwZgySj5Tk1+as+v1PKe3+uxPlOm25PLheJK52mGWe4ggGZx0CY2VOkD/g7
kRRs+w+CFXPV62/zSgDLMlhCfnK8PoYs7uQoybm6zgECZc+2MPOAeHKN/MWPOdZv
zUipIcQQ9mhl/E2NmncLiSefZbZx6hU7wmfzAywQSvlRyU2PRS5p/vckKkID36xU
xI/v/JR6oudBkQYpqrcz4ulzc4bbrX4BY8oueT1rzPWgIBNsZUPe1+p7oOTzJ7Ze
OFBUTsB3DtcPOGVbMD3RBmiqbNtWQzqfjyyd01f2D4Tz4yGN+XWp7oqVzxvoe+Ad
TgPC3FYVJ+va481hDCdSAZGctola7rWZVQBxPON6TBQuzw32bSy1ySYh6yLgRphm
nRdTnmEBdiwBryXhnPe7XGHaRyubqhJFBG3FAip+rLg66aXmfPzWEfLybKWIWv1D
zpbobssIK9xGndf//0CmrY4+9en1RjIcjOU+EH09GqWhyU+YGGZvZJjt/PWu2V4J
o3CR/fouKoJ1ibkBbopOW4UfYREbu/fYnkiTcddfIGdzvUQFv+bzbnNTW+A575k6
d+gLAI1PYQPAhYds4JpjBDSGVM/1zdFGy1niNfxfjE9Ohk8Ljo2Aole3nVbOdMAd
3Ff2EvfUuK/lah5MUmS2TCN2C8K9yS/Skg9eeHVIRza8KmFKxreoMuvZ5dSIC6nY
eCp1J0TZibYIgOME002JcdBjFXUZv+Dng+Fh1Uc4kHGCybU1GgEJyKb8jFeH6f9/
ND9d6bDGbnlWz6sZd5y4+bgeUWVFfbgUKo4Ocp7T05a+o3ucao1MW41y/G/gkhqk
SS3imPjwFKowe5ppsjzoPeOEoCIeTheWfk6+H7EELoBK/nk5z2LT6DEpFSromSVz
VCBsoXWOLNUdiyBvsc/Xwdx5h6P5EJMsKoO2PCDqLYzNDj2EqCkZk1KjbKOk0h3q
KU+VCSc1NUyEX5277oaXNTi1KBE464riTa4vbWHP61LfLURcD+/JIxgUQBNU2CIf
LVq0nEquGmS7YxT9j0EZMh8veU5zctoOyEhnGYctRqPYYjqbHaY0S0+03wSxOMa6
Ztt6POHexKc693xCNflC4zWulCzNnHz+oDervdtRZ4w6Onjw7UIuk+Av7Lwbl3Gg
jZXwqLqJ4qgo8/6Zx0d+d/WSO45xsklZbPtQ7/EGoBa/DHvNTtO2OSpYwvKIEEcq
qleSNhSmoxaAz0R/b8ni/C3JAQ+PRQLs/sQ7XQR9YNEX4cCmIK3a7z8DdMNPloEy
S8a6wz1LUgdB5Y7Pfc1vxWCuL6HpiqWzXJeA7lWAcm8k4bamwg8SEvnJXRXTz326
p8KzSPUDsSlzWnn1jhgqbgCs1tOLYURfu+XBoKjtx1mAqGo+VVFYlyI1CLwgpzHW
jSfLr4YDLGh6/7HmI3KbHKs/WlopyFY620TvLjC21AQtaFR1Z0mm2Jfv95O3T9oO
0Ad+38JccBNgVYS7Fs1Pqi3WAJd6fiEt1JvUV9VIfSuAOtMiXWadNnnNZ0OSqobf
XsIaeVfu+deWttm9FivPdOAYTT4Nny5CGaXny7raS30JklofGHx1bu1le4fwqGci
7fL+eGGn0IcNcp7HQeLXuUq5t/1bq7sUXOp9Ul0c85dDF1hsUc51wEBBXawgn3q2
4IoG4Yj9aWJfZwVHscu1V/nvqsfqgniuXeGJ3RuWtihV8BUgR/CEJjjUgbOp9x13
mTLP8Zh4WHajQ0GCdJsEe8l1uhHGWz2KtJZoKy839F+vGRFaphtqXPVkSz7vvYXV
bco3lL+U+LVo1/yDB8FKG/mBC6tXetV35ufVT7sl+NT0qFYAYg6bdrEun+tVnCHg
3I0u9d3K2IeNi/zQE2JJo+w8+PcyzcOkeWu2PU/91+iiChU0GKW0B4oSf17NCEuY
eHMDpGAmUEPxEqssmsdfwZHpacE5c0TkTrXaK7wNK8CP1koQIJIz+sEW/CC1f+nn
SD9iMrOjYjfkDCCFd0ALe7hJsoBlUplklDbZXyIbyJwP9BBWQbpsZuVZkJz/PD5M
r0ZmhcGGmWzWLHJyVKQubXQd8yNt3VpwQexHHjhza41vH3Xt735clLJtZex/7NEj
bu53MMw18aXWy/pMRvDPv2iv+jORn6Pgujy8Fquy1CWyvUG9sUxqUW0JH4Qy3TWf
C7tBgKVfqtFPX3BQCHpg0Q==
`pragma protect end_protected
