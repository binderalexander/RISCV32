-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- VENDOR "Altera"
-- PROGRAM "Quartus Prime"
-- VERSION "Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition"

-- DATE "05/17/2020 18:22:12"

-- 
-- Device: Altera 5CSEMA5F31C6 Package FBGA896
-- 

-- 
-- This VHDL file should be used for ModelSim (VHDL) only
-- 

LIBRARY ALTERA;
LIBRARY ALTERA_LNSIM;
LIBRARY CYCLONEV;
LIBRARY IEEE;
USE ALTERA.ALTERA_PRIMITIVES_COMPONENTS.ALL;
USE ALTERA_LNSIM.ALTERA_LNSIM_COMPONENTS.ALL;
USE CYCLONEV.CYCLONEV_COMPONENTS.ALL;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY 	Core IS
    PORT (
	csi_clk : IN std_logic;
	rsi_reset_n : IN std_logic;
	avm_i_address : OUT std_logic_vector(31 DOWNTO 0);
	avm_i_read : OUT std_logic;
	avm_i_readdata : IN std_logic_vector(31 DOWNTO 0);
	avm_i_waitrequest : IN std_logic;
	avm_d_address : OUT std_logic_vector(31 DOWNTO 0);
	avm_d_byteenable : OUT std_logic_vector(3 DOWNTO 0);
	avm_d_write : OUT std_logic;
	avm_d_writedata : OUT std_logic_vector(31 DOWNTO 0);
	avm_d_read : OUT std_logic;
	avm_d_readdata : IN std_logic_vector(31 DOWNTO 0);
	avm_d_waitrequest : IN std_logic
	);
END Core;

-- Design Ports Information
-- avm_i_address[0]	=>  Location: PIN_H15,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[1]	=>  Location: PIN_AF13,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[2]	=>  Location: PIN_W24,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[3]	=>  Location: PIN_AD26,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[4]	=>  Location: PIN_AF29,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[5]	=>  Location: PIN_AE27,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[6]	=>  Location: PIN_V23,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[7]	=>  Location: PIN_AF28,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[8]	=>  Location: PIN_Y23,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[9]	=>  Location: PIN_AC23,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[10]	=>  Location: PIN_AE26,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[11]	=>  Location: PIN_Y21,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[12]	=>  Location: PIN_W21,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[13]	=>  Location: PIN_AE28,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[14]	=>  Location: PIN_AJ29,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[15]	=>  Location: PIN_AH29,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[16]	=>  Location: PIN_AG27,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[17]	=>  Location: PIN_AJ20,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[18]	=>  Location: PIN_AF21,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[19]	=>  Location: PIN_W20,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[20]	=>  Location: PIN_W22,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[21]	=>  Location: PIN_AF19,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[22]	=>  Location: PIN_AD21,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[23]	=>  Location: PIN_AH28,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[24]	=>  Location: PIN_AC25,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[25]	=>  Location: PIN_AD20,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[26]	=>  Location: PIN_AF20,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[27]	=>  Location: PIN_AK28,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[28]	=>  Location: PIN_AK24,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[29]	=>  Location: PIN_AE24,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[30]	=>  Location: PIN_AF14,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_address[31]	=>  Location: PIN_AG13,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_read	=>  Location: PIN_AJ17,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_waitrequest	=>  Location: PIN_E3,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[0]	=>  Location: PIN_AH30,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[1]	=>  Location: PIN_AG28,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[2]	=>  Location: PIN_AA24,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[3]	=>  Location: PIN_AB22,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[4]	=>  Location: PIN_A11,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[5]	=>  Location: PIN_AD27,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[6]	=>  Location: PIN_AB23,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[7]	=>  Location: PIN_AA25,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[8]	=>  Location: PIN_C13,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[9]	=>  Location: PIN_AH7,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[10]	=>  Location: PIN_AC29,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[11]	=>  Location: PIN_AC27,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[12]	=>  Location: PIN_A10,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[13]	=>  Location: PIN_AF30,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[14]	=>  Location: PIN_AK6,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[15]	=>  Location: PIN_AB30,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[16]	=>  Location: PIN_AH12,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[17]	=>  Location: PIN_AH14,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[18]	=>  Location: PIN_AH13,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[19]	=>  Location: PIN_AF26,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[20]	=>  Location: PIN_V25,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[21]	=>  Location: PIN_AK18,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[22]	=>  Location: PIN_AJ19,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[23]	=>  Location: PIN_AC22,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[24]	=>  Location: PIN_AF25,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[25]	=>  Location: PIN_AB26,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[26]	=>  Location: PIN_AJ5,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[27]	=>  Location: PIN_AC28,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[28]	=>  Location: PIN_AG12,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[29]	=>  Location: PIN_AA21,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[30]	=>  Location: PIN_D11,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_address[31]	=>  Location: PIN_B13,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_byteenable[0]	=>  Location: PIN_AD24,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_byteenable[1]	=>  Location: PIN_AG17,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_byteenable[2]	=>  Location: PIN_AK8,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_byteenable[3]	=>  Location: PIN_AB15,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_write	=>  Location: PIN_AH8,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[0]	=>  Location: PIN_AH17,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[1]	=>  Location: PIN_AG21,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[2]	=>  Location: PIN_AH20,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[3]	=>  Location: PIN_AJ9,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[4]	=>  Location: PIN_AK7,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[5]	=>  Location: PIN_AJ16,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[6]	=>  Location: PIN_AK12,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[7]	=>  Location: PIN_AK9,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[8]	=>  Location: PIN_W17,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[9]	=>  Location: PIN_W16,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[10]	=>  Location: PIN_AA16,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[11]	=>  Location: PIN_B12,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[12]	=>  Location: PIN_V16,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[13]	=>  Location: PIN_AF18,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[14]	=>  Location: PIN_AE16,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[15]	=>  Location: PIN_AB17,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[16]	=>  Location: PIN_AG2,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[17]	=>  Location: PIN_AH15,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[18]	=>  Location: PIN_AG15,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[19]	=>  Location: PIN_AC14,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[20]	=>  Location: PIN_AK14,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[21]	=>  Location: PIN_AE17,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[22]	=>  Location: PIN_W15,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[23]	=>  Location: PIN_AF16,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[24]	=>  Location: PIN_AG16,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[25]	=>  Location: PIN_AD25,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[26]	=>  Location: PIN_AG30,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[27]	=>  Location: PIN_AJ14,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[28]	=>  Location: PIN_AJ12,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[29]	=>  Location: PIN_A13,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[30]	=>  Location: PIN_Y16,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_writedata[31]	=>  Location: PIN_G15,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_read	=>  Location: PIN_AJ11,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_waitrequest	=>  Location: PIN_B8,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- csi_clk	=>  Location: PIN_Y27,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- rsi_reset_n	=>  Location: PIN_AA26,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[21]	=>  Location: PIN_AK27,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[22]	=>  Location: PIN_W19,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[20]	=>  Location: PIN_AE23,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[14]	=>  Location: PIN_AH22,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[12]	=>  Location: PIN_AG22,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[13]	=>  Location: PIN_AE19,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[15]	=>  Location: PIN_AJ22,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[0]	=>  Location: PIN_Y18,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[27]	=>  Location: PIN_AH25,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[29]	=>  Location: PIN_AK26,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[28]	=>  Location: PIN_AJ26,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[30]	=>  Location: PIN_AC20,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[26]	=>  Location: PIN_AD19,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[25]	=>  Location: PIN_AE22,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[24]	=>  Location: PIN_AG25,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[2]	=>  Location: PIN_AK29,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[3]	=>  Location: PIN_AJ27,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[4]	=>  Location: PIN_AJ25,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[5]	=>  Location: PIN_V18,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[6]	=>  Location: PIN_AJ24,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[7]	=>  Location: PIN_AF24,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[1]	=>  Location: PIN_AF23,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[9]	=>  Location: PIN_AC18,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[23]	=>  Location: PIN_AH24,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[8]	=>  Location: PIN_AD17,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[10]	=>  Location: PIN_AG23,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[11]	=>  Location: PIN_AE18,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[31]	=>  Location: PIN_AA19,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[16]	=>  Location: PIN_AK22,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[18]	=>  Location: PIN_AK21,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[17]	=>  Location: PIN_AA18,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_i_readdata[19]	=>  Location: PIN_Y17,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[0]	=>  Location: PIN_AK23,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[31]	=>  Location: PIN_AG26,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[23]	=>  Location: PIN_AA20,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[16]	=>  Location: PIN_AJ21,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[24]	=>  Location: PIN_AH23,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[1]	=>  Location: PIN_AB21,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[17]	=>  Location: PIN_AF15,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[25]	=>  Location: PIN_AA28,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[2]	=>  Location: PIN_F14,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[18]	=>  Location: PIN_AH18,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[26]	=>  Location: PIN_Y24,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[3]	=>  Location: PIN_AH27,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[19]	=>  Location: PIN_A8,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[27]	=>  Location: PIN_W25,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[4]	=>  Location: PIN_AH10,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[20]	=>  Location: PIN_AG20,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[28]	=>  Location: PIN_AB28,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[5]	=>  Location: PIN_AB13,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[21]	=>  Location: PIN_AA15,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[29]	=>  Location: PIN_AB25,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[6]	=>  Location: PIN_AK16,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[22]	=>  Location: PIN_AK19,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[30]	=>  Location: PIN_C12,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[7]	=>  Location: PIN_AE13,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[8]	=>  Location: PIN_V17,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[9]	=>  Location: PIN_AH19,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[10]	=>  Location: PIN_AJ10,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[11]	=>  Location: PIN_AG18,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[12]	=>  Location: PIN_AK13,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[13]	=>  Location: PIN_Y19,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[14]	=>  Location: PIN_AK11,	 I/O Standard: 2.5 V,	 Current Strength: Default
-- avm_d_readdata[15]	=>  Location: PIN_AA14,	 I/O Standard: 2.5 V,	 Current Strength: Default


ARCHITECTURE structure OF Core IS
SIGNAL gnd : std_logic := '0';
SIGNAL vcc : std_logic := '1';
SIGNAL unknown : std_logic := 'X';
SIGNAL devoe : std_logic := '1';
SIGNAL devclrn : std_logic := '1';
SIGNAL devpor : std_logic := '1';
SIGNAL ww_devoe : std_logic;
SIGNAL ww_devclrn : std_logic;
SIGNAL ww_devpor : std_logic;
SIGNAL ww_csi_clk : std_logic;
SIGNAL ww_rsi_reset_n : std_logic;
SIGNAL ww_avm_i_address : std_logic_vector(31 DOWNTO 0);
SIGNAL ww_avm_i_read : std_logic;
SIGNAL ww_avm_i_readdata : std_logic_vector(31 DOWNTO 0);
SIGNAL ww_avm_i_waitrequest : std_logic;
SIGNAL ww_avm_d_address : std_logic_vector(31 DOWNTO 0);
SIGNAL ww_avm_d_byteenable : std_logic_vector(3 DOWNTO 0);
SIGNAL ww_avm_d_write : std_logic;
SIGNAL ww_avm_d_writedata : std_logic_vector(31 DOWNTO 0);
SIGNAL ww_avm_d_read : std_logic;
SIGNAL ww_avm_d_readdata : std_logic_vector(31 DOWNTO 0);
SIGNAL ww_avm_d_waitrequest : std_logic;
SIGNAL \avm_i_waitrequest~input_o\ : std_logic;
SIGNAL \avm_d_waitrequest~input_o\ : std_logic;
SIGNAL \csi_clk~input_o\ : std_logic;
SIGNAL \csi_clk~inputCLKENA0_outclk\ : std_logic;
SIGNAL \avm_i_readdata[31]~input_o\ : std_logic;
SIGNAL \rsi_reset_n~input_o\ : std_logic;
SIGNAL \rsi_reset_n~inputCLKENA0_outclk\ : std_logic;
SIGNAL \avm_i_readdata[26]~input_o\ : std_logic;
SIGNAL \avm_i_readdata[28]~input_o\ : std_logic;
SIGNAL \avm_i_readdata[30]~input_o\ : std_logic;
SIGNAL \avm_i_readdata[29]~input_o\ : std_logic;
SIGNAL \avm_i_readdata[12]~input_o\ : std_logic;
SIGNAL \Mux154~1_combout\ : std_logic;
SIGNAL \avm_i_readdata[27]~input_o\ : std_logic;
SIGNAL \avm_i_readdata[24]~input_o\ : std_logic;
SIGNAL \avm_i_readdata[25]~input_o\ : std_logic;
SIGNAL \Equal4~1_combout\ : std_logic;
SIGNAL \Mux34~0_combout\ : std_logic;
SIGNAL \avm_i_readdata[22]~input_o\ : std_logic;
SIGNAL \avm_i_readdata[21]~input_o\ : std_logic;
SIGNAL \avm_i_readdata[20]~input_o\ : std_logic;
SIGNAL \Mux0~0_combout\ : std_logic;
SIGNAL \Mux11~0_combout\ : std_logic;
SIGNAL \NxR~12_combout\ : std_logic;
SIGNAL \R.ctrlState.Calc~q\ : std_logic;
SIGNAL \Mux53~0_combout\ : std_logic;
SIGNAL \R.ctrlState.DataAccess0~DUPLICATE_q\ : std_logic;
SIGNAL \Mux50~0_combout\ : std_logic;
SIGNAL \NxR~13_combout\ : std_logic;
SIGNAL \R.ctrlState.DataAccess0~q\ : std_logic;
SIGNAL \Mux18~0_combout\ : std_logic;
SIGNAL \Mux53~1_combout\ : std_logic;
SIGNAL \Mux53~2_combout\ : std_logic;
SIGNAL \avm_i_readdata[3]~input_o\ : std_logic;
SIGNAL \avm_i_readdata[5]~input_o\ : std_logic;
SIGNAL \avm_i_readdata[6]~input_o\ : std_logic;
SIGNAL \avm_i_readdata[4]~input_o\ : std_logic;
SIGNAL \avm_i_readdata[7]~input_o\ : std_logic;
SIGNAL \Equal2~0_combout\ : std_logic;
SIGNAL \avm_i_readdata[2]~input_o\ : std_logic;
SIGNAL \avm_i_readdata[14]~input_o\ : std_logic;
SIGNAL \avm_i_readdata[15]~input_o\ : std_logic;
SIGNAL \avm_i_readdata[1]~input_o\ : std_logic;
SIGNAL \avm_i_readdata[0]~input_o\ : std_logic;
SIGNAL \Equal2~1_combout\ : std_logic;
SIGNAL \avm_i_readdata[13]~input_o\ : std_logic;
SIGNAL \Equal2~2_combout\ : std_logic;
SIGNAL \NxR~20_combout\ : std_logic;
SIGNAL \R.ctrlState.Trap~q\ : std_logic;
SIGNAL \NxR~18_combout\ : std_logic;
SIGNAL \R.ctrlState.CheckJump~q\ : std_logic;
SIGNAL \Mux154~0_combout\ : std_logic;
SIGNAL \NxR~4_combout\ : std_logic;
SIGNAL \Mux12~0_combout\ : std_logic;
SIGNAL \NxR~14_combout\ : std_logic;
SIGNAL \R.ctrlState.Wait0~q\ : std_logic;
SIGNAL \NxR~0_combout\ : std_logic;
SIGNAL \NxR~1_combout\ : std_logic;
SIGNAL \R.ctrlState.Wait1~q\ : std_logic;
SIGNAL \vAluSrc1~0_combout\ : std_logic;
SIGNAL \Mux123~0_combout\ : std_logic;
SIGNAL \NxR~2_combout\ : std_logic;
SIGNAL \NxR~15_combout\ : std_logic;
SIGNAL \NxR~16_combout\ : std_logic;
SIGNAL \R.ctrlState.DataAccess1~q\ : std_logic;
SIGNAL \NxR~3_combout\ : std_logic;
SIGNAL \R.ctrlState.WriteReg~q\ : std_logic;
SIGNAL \Comb~0_combout\ : std_logic;
SIGNAL \NxR~17_combout\ : std_logic;
SIGNAL \R.ctrlState.Fetch~q\ : std_logic;
SIGNAL \R.ctrlState.ReadReg~q\ : std_logic;
SIGNAL \vAluSrc2~0_combout\ : std_logic;
SIGNAL \vAluSrc2~1_combout\ : std_logic;
SIGNAL \~GND~combout\ : std_logic;
SIGNAL \R.memToReg~q\ : std_logic;
SIGNAL \avm_d_readdata[24]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[0]~0_combout\ : std_logic;
SIGNAL \NxR~5_combout\ : std_logic;
SIGNAL \R.aluCalc~q\ : std_logic;
SIGNAL \Mux124~0_combout\ : std_logic;
SIGNAL \Mux123~1_combout\ : std_logic;
SIGNAL \Mux131~0_combout\ : std_logic;
SIGNAL \Comb~1_combout\ : std_logic;
SIGNAL \Mux18~1_combout\ : std_logic;
SIGNAL \Mux18~2_combout\ : std_logic;
SIGNAL \R.aluOp.ALUOpSub~q\ : std_logic;
SIGNAL \Mux17~0_combout\ : std_logic;
SIGNAL \Mux17~1_combout\ : std_logic;
SIGNAL \R.aluOp.ALUOpAdd_OTERM365\ : std_logic;
SIGNAL \R.aluOp.ALUOpAdd~q\ : std_logic;
SIGNAL \vAluSrc1~2_combout\ : std_logic;
SIGNAL \vAluSrc1~1_combout\ : std_logic;
SIGNAL \avm_i_readdata[10]~input_o\ : std_logic;
SIGNAL \avm_i_readdata[11]~input_o\ : std_logic;
SIGNAL \avm_i_readdata[19]~input_o\ : std_logic;
SIGNAL \avm_i_readdata[18]~input_o\ : std_logic;
SIGNAL \avm_i_readdata[17]~input_o\ : std_logic;
SIGNAL \avm_i_readdata[16]~input_o\ : std_logic;
SIGNAL \Mux31~0_combout\ : std_logic;
SIGNAL \NxR~19_combout\ : std_logic;
SIGNAL \R.csrRead~q\ : std_logic;
SIGNAL \R.regWriteEn~1_combout\ : std_logic;
SIGNAL \R.regWriteEn~0_combout\ : std_logic;
SIGNAL \R.regWriteEn~2_combout\ : std_logic;
SIGNAL \R.regWriteEn~q\ : std_logic;
SIGNAL \Decoder0~11_combout\ : std_logic;
SIGNAL \RegFile[21][23]~q\ : std_logic;
SIGNAL \Decoder0~12_combout\ : std_logic;
SIGNAL \RegFile[23][23]~q\ : std_logic;
SIGNAL \RegFile[22][23]~feeder_combout\ : std_logic;
SIGNAL \Decoder0~14_combout\ : std_logic;
SIGNAL \RegFile[22][23]~q\ : std_logic;
SIGNAL \avm_i_readdata[9]~input_o\ : std_logic;
SIGNAL \avm_i_readdata[8]~input_o\ : std_logic;
SIGNAL \Decoder0~24_combout\ : std_logic;
SIGNAL \RegFile[19][23]~q\ : std_logic;
SIGNAL \Decoder0~23_combout\ : std_logic;
SIGNAL \RegFile[17][23]~q\ : std_logic;
SIGNAL \Decoder0~26_combout\ : std_logic;
SIGNAL \RegFile[18][23]~q\ : std_logic;
SIGNAL \avm_i_readdata[23]~input_o\ : std_logic;
SIGNAL \RegFile[16][23]~feeder_combout\ : std_logic;
SIGNAL \Decoder0~25_combout\ : std_logic;
SIGNAL \RegFile[16][23]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux67~18_combout\ : std_logic;
SIGNAL \RegFile[20][23]~feeder_combout\ : std_logic;
SIGNAL \Decoder0~13_combout\ : std_logic;
SIGNAL \RegFile[20][23]~q\ : std_logic;
SIGNAL \Mux67~5_combout\ : std_logic;
SIGNAL \Decoder0~10_combout\ : std_logic;
SIGNAL \RegFile[14][23]~q\ : std_logic;
SIGNAL \Decoder0~7_combout\ : std_logic;
SIGNAL \RegFile[13][23]~q\ : std_logic;
SIGNAL \Decoder0~20_combout\ : std_logic;
SIGNAL \RegFile[11][23]~q\ : std_logic;
SIGNAL \Decoder0~22_combout\ : std_logic;
SIGNAL \RegFile[10][23]~q\ : std_logic;
SIGNAL \Decoder0~19_combout\ : std_logic;
SIGNAL \RegFile[9][23]~q\ : std_logic;
SIGNAL \RegFile[8][23]~feeder_combout\ : std_logic;
SIGNAL \Decoder0~21_combout\ : std_logic;
SIGNAL \RegFile[8][23]~q\ : std_logic;
SIGNAL \Mux67~14_combout\ : std_logic;
SIGNAL \Decoder0~9_combout\ : std_logic;
SIGNAL \RegFile[12][23]~q\ : std_logic;
SIGNAL \Mux67~1_combout\ : std_logic;
SIGNAL \Decoder0~6_combout\ : std_logic;
SIGNAL \RegFile[3][23]~q\ : std_logic;
SIGNAL \Decoder0~4_combout\ : std_logic;
SIGNAL \RegFile[2][23]~q\ : std_logic;
SIGNAL \Decoder0~2_combout\ : std_logic;
SIGNAL \RegFile[6][23]~q\ : std_logic;
SIGNAL \Decoder0~0_combout\ : std_logic;
SIGNAL \RegFile[4][23]~q\ : std_logic;
SIGNAL \RegFile[5][23]~feeder_combout\ : std_logic;
SIGNAL \Decoder0~1_combout\ : std_logic;
SIGNAL \RegFile[5][23]~q\ : std_logic;
SIGNAL \Decoder0~3_combout\ : std_logic;
SIGNAL \RegFile[7][23]~q\ : std_logic;
SIGNAL \Mux67~0_combout\ : std_logic;
SIGNAL \RegFile[1][23]~feeder_combout\ : std_logic;
SIGNAL \Decoder0~5_combout\ : std_logic;
SIGNAL \RegFile[1][23]~q\ : std_logic;
SIGNAL \Mux67~26_combout\ : std_logic;
SIGNAL \Decoder0~16_combout\ : std_logic;
SIGNAL \RegFile[31][23]~q\ : std_logic;
SIGNAL \Decoder0~15_combout\ : std_logic;
SIGNAL \RegFile[29][23]~q\ : std_logic;
SIGNAL \RegFile[30][23]~feeder_combout\ : std_logic;
SIGNAL \Decoder0~18_combout\ : std_logic;
SIGNAL \RegFile[30][23]~q\ : std_logic;
SIGNAL \Decoder0~28_combout\ : std_logic;
SIGNAL \RegFile[27][23]~q\ : std_logic;
SIGNAL \Decoder0~30_combout\ : std_logic;
SIGNAL \RegFile[26][23]~q\ : std_logic;
SIGNAL \Decoder0~27_combout\ : std_logic;
SIGNAL \RegFile[25][23]~q\ : std_logic;
SIGNAL \RegFile[24][23]~feeder_combout\ : std_logic;
SIGNAL \Decoder0~29_combout\ : std_logic;
SIGNAL \RegFile[24][23]~q\ : std_logic;
SIGNAL \Mux67~22_combout\ : std_logic;
SIGNAL \RegFile[28][23]~feeder_combout\ : std_logic;
SIGNAL \Decoder0~17_combout\ : std_logic;
SIGNAL \RegFile[28][23]~q\ : std_logic;
SIGNAL \Mux67~9_combout\ : std_logic;
SIGNAL \Mux67~13_combout\ : std_logic;
SIGNAL \Mux231~0_combout\ : std_logic;
SIGNAL \Mux132~0_combout\ : std_logic;
SIGNAL \Equal4~0_combout\ : std_logic;
SIGNAL \Equal4~2_combout\ : std_logic;
SIGNAL \RegFile[21][22]~q\ : std_logic;
SIGNAL \RegFile[23][22]~q\ : std_logic;
SIGNAL \RegFile[22][22]~q\ : std_logic;
SIGNAL \RegFile[17][22]~q\ : std_logic;
SIGNAL \RegFile[19][22]~q\ : std_logic;
SIGNAL \RegFile[18][22]~feeder_combout\ : std_logic;
SIGNAL \RegFile[18][22]~q\ : std_logic;
SIGNAL \RegFile[16][22]~feeder_combout\ : std_logic;
SIGNAL \RegFile[16][22]~q\ : std_logic;
SIGNAL \Mux68~18_combout\ : std_logic;
SIGNAL \RegFile[20][22]~q\ : std_logic;
SIGNAL \Mux68~5_combout\ : std_logic;
SIGNAL \RegFile[30][22]~q\ : std_logic;
SIGNAL \RegFile[29][22]~q\ : std_logic;
SIGNAL \RegFile[27][22]~q\ : std_logic;
SIGNAL \RegFile[25][22]~q\ : std_logic;
SIGNAL \RegFile[26][22]~feeder_combout\ : std_logic;
SIGNAL \RegFile[26][22]~q\ : std_logic;
SIGNAL \RegFile[24][22]~feeder_combout\ : std_logic;
SIGNAL \RegFile[24][22]~q\ : std_logic;
SIGNAL \Mux68~22_combout\ : std_logic;
SIGNAL \RegFile[28][22]~q\ : std_logic;
SIGNAL \Mux68~9_combout\ : std_logic;
SIGNAL \RegFile[3][22]~q\ : std_logic;
SIGNAL \RegFile[2][22]~q\ : std_logic;
SIGNAL \RegFile[4][22]~feeder_combout\ : std_logic;
SIGNAL \RegFile[4][22]~q\ : std_logic;
SIGNAL \RegFile[5][22]~q\ : std_logic;
SIGNAL \RegFile[6][22]~q\ : std_logic;
SIGNAL \RegFile[7][22]~q\ : std_logic;
SIGNAL \Mux68~0_combout\ : std_logic;
SIGNAL \RegFile[1][22]~feeder_combout\ : std_logic;
SIGNAL \RegFile[1][22]~q\ : std_logic;
SIGNAL \Mux68~26_combout\ : std_logic;
SIGNAL \RegFile[13][22]~q\ : std_logic;
SIGNAL \RegFile[14][22]~feeder_combout\ : std_logic;
SIGNAL \RegFile[14][22]~q\ : std_logic;
SIGNAL \Decoder0~8_combout\ : std_logic;
SIGNAL \RegFile[15][22]~q\ : std_logic;
SIGNAL \RegFile[11][22]~q\ : std_logic;
SIGNAL \RegFile[10][22]~feeder_combout\ : std_logic;
SIGNAL \RegFile[10][22]~q\ : std_logic;
SIGNAL \RegFile[9][22]~q\ : std_logic;
SIGNAL \RegFile[8][22]~q\ : std_logic;
SIGNAL \Mux68~14_combout\ : std_logic;
SIGNAL \RegFile[12][22]~feeder_combout\ : std_logic;
SIGNAL \RegFile[12][22]~q\ : std_logic;
SIGNAL \Mux68~1_combout\ : std_logic;
SIGNAL \Mux68~13_combout\ : std_logic;
SIGNAL \Mux232~0_combout\ : std_logic;
SIGNAL \R.aluOp.ALUOpSLL~q\ : std_logic;
SIGNAL \Mux26~0_combout\ : std_logic;
SIGNAL \Mux162~0_combout\ : std_logic;
SIGNAL \Mux24~0_combout\ : std_logic;
SIGNAL \Mux24~1_combout\ : std_logic;
SIGNAL \R.aluOp.ALUOpSLL_OTERM359\ : std_logic;
SIGNAL \Mux150~0_combout\ : std_logic;
SIGNAL \R.aluOp.ALUOpSRL~q\ : std_logic;
SIGNAL \Mux21~0_combout\ : std_logic;
SIGNAL \Mux25~0_combout\ : std_logic;
SIGNAL \Mux25~1_combout\ : std_logic;
SIGNAL \R.aluOp.ALUOpSRL_OTERM361\ : std_logic;
SIGNAL \Selector31~7_combout\ : std_logic;
SIGNAL \Selector31~7_OTERM383\ : std_logic;
SIGNAL \Selector31~0_OTERM349\ : std_logic;
SIGNAL \R.aluOp.ALUOpSRA_OTERM363\ : std_logic;
SIGNAL \R.aluOp.ALUOpSRA~q\ : std_logic;
SIGNAL \Mux26~1_combout\ : std_logic;
SIGNAL \Mux26~2_combout\ : std_logic;
SIGNAL \Selector31~0_NEW_REG348_OTERM569\ : std_logic;
SIGNAL \Selector31~5_combout\ : std_logic;
SIGNAL \Selector31~5_OTERM599\ : std_logic;
SIGNAL \Mux152~0_combout\ : std_logic;
SIGNAL \Selector31~6_combout\ : std_logic;
SIGNAL \Selector31~6_OTERM381\ : std_logic;
SIGNAL \Mux127~0_combout\ : std_logic;
SIGNAL \Mux123~3_combout\ : std_logic;
SIGNAL \RegFile[2][21]~q\ : std_logic;
SIGNAL \RegFile[5][21]~q\ : std_logic;
SIGNAL \RegFile[6][21]~feeder_combout\ : std_logic;
SIGNAL \RegFile[6][21]~q\ : std_logic;
SIGNAL \RegFile[4][21]~feeder_combout\ : std_logic;
SIGNAL \RegFile[4][21]~q\ : std_logic;
SIGNAL \RegFile[7][21]~q\ : std_logic;
SIGNAL \Mux69~0_combout\ : std_logic;
SIGNAL \RegFile[1][21]~feeder_combout\ : std_logic;
SIGNAL \RegFile[1][21]~q\ : std_logic;
SIGNAL \Mux69~26_combout\ : std_logic;
SIGNAL \RegFile[13][21]~q\ : std_logic;
SIGNAL \RegFile[14][21]~feeder_combout\ : std_logic;
SIGNAL \RegFile[14][21]~q\ : std_logic;
SIGNAL \RegFile[15][21]~q\ : std_logic;
SIGNAL \RegFile[9][21]~q\ : std_logic;
SIGNAL \RegFile[11][21]~q\ : std_logic;
SIGNAL \RegFile[10][21]~feeder_combout\ : std_logic;
SIGNAL \RegFile[10][21]~q\ : std_logic;
SIGNAL \RegFile[8][21]~feeder_combout\ : std_logic;
SIGNAL \RegFile[8][21]~q\ : std_logic;
SIGNAL \Mux69~14_combout\ : std_logic;
SIGNAL \RegFile[12][21]~q\ : std_logic;
SIGNAL \Mux69~1_combout\ : std_logic;
SIGNAL \RegFile[31][21]~q\ : std_logic;
SIGNAL \RegFile[29][21]~q\ : std_logic;
SIGNAL \RegFile[30][21]~q\ : std_logic;
SIGNAL \RegFile[27][21]~q\ : std_logic;
SIGNAL \RegFile[25][21]~q\ : std_logic;
SIGNAL \RegFile[26][21]~feeder_combout\ : std_logic;
SIGNAL \RegFile[26][21]~q\ : std_logic;
SIGNAL \RegFile[24][21]~feeder_combout\ : std_logic;
SIGNAL \RegFile[24][21]~q\ : std_logic;
SIGNAL \Mux69~22_combout\ : std_logic;
SIGNAL \RegFile[28][21]~feeder_combout\ : std_logic;
SIGNAL \RegFile[28][21]~q\ : std_logic;
SIGNAL \Mux69~9_combout\ : std_logic;
SIGNAL \RegFile[23][21]~q\ : std_logic;
SIGNAL \RegFile[22][21]~q\ : std_logic;
SIGNAL \RegFile[21][21]~q\ : std_logic;
SIGNAL \RegFile[19][21]~q\ : std_logic;
SIGNAL \RegFile[18][21]~feeder_combout\ : std_logic;
SIGNAL \RegFile[18][21]~q\ : std_logic;
SIGNAL \RegFile[17][21]~q\ : std_logic;
SIGNAL \RegFile[16][21]~feeder_combout\ : std_logic;
SIGNAL \RegFile[16][21]~q\ : std_logic;
SIGNAL \Mux69~18_combout\ : std_logic;
SIGNAL \RegFile[20][21]~feeder_combout\ : std_logic;
SIGNAL \RegFile[20][21]~q\ : std_logic;
SIGNAL \Mux69~5_combout\ : std_logic;
SIGNAL \Mux69~13_combout\ : std_logic;
SIGNAL \Mux233~0_combout\ : std_logic;
SIGNAL \Mux153~0_combout\ : std_logic;
SIGNAL \Mux222~0_combout\ : std_logic;
SIGNAL \avm_d_readdata[25]~input_o\ : std_logic;
SIGNAL \Add2~1_OTERM735_OTERM839\ : std_logic;
SIGNAL \RegFile[31][0]~q\ : std_logic;
SIGNAL \RegFile[30][0]~q\ : std_logic;
SIGNAL \RegFile[29][0]~q\ : std_logic;
SIGNAL \RegFile[25][0]~q\ : std_logic;
SIGNAL \RegFile[26][0]~q\ : std_logic;
SIGNAL \RegFile[27][0]~q\ : std_logic;
SIGNAL \RegFile[24][0]~feeder_combout\ : std_logic;
SIGNAL \RegFile[24][0]~q\ : std_logic;
SIGNAL \Mux90~22_combout\ : std_logic;
SIGNAL \RegFile[28][0]~feeder_combout\ : std_logic;
SIGNAL \RegFile[28][0]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux90~9_combout\ : std_logic;
SIGNAL \RegFile[2][0]~q\ : std_logic;
SIGNAL \RegFile[4][0]~feeder_combout\ : std_logic;
SIGNAL \RegFile[4][0]~q\ : std_logic;
SIGNAL \RegFile[6][0]~feeder_combout\ : std_logic;
SIGNAL \RegFile[6][0]~q\ : std_logic;
SIGNAL \RegFile[5][0]~feeder_combout\ : std_logic;
SIGNAL \RegFile[5][0]~q\ : std_logic;
SIGNAL \RegFile[7][0]~feeder_combout\ : std_logic;
SIGNAL \RegFile[7][0]~q\ : std_logic;
SIGNAL \Mux90~0_combout\ : std_logic;
SIGNAL \RegFile[1][0]~feeder_combout\ : std_logic;
SIGNAL \RegFile[1][0]~q\ : std_logic;
SIGNAL \Mux90~26_combout\ : std_logic;
SIGNAL \RegFile[13][0]~q\ : std_logic;
SIGNAL \RegFile[14][0]~feeder_combout\ : std_logic;
SIGNAL \RegFile[14][0]~q\ : std_logic;
SIGNAL \RegFile[15][0]~q\ : std_logic;
SIGNAL \RegFile[11][0]~q\ : std_logic;
SIGNAL \RegFile[9][0]~feeder_combout\ : std_logic;
SIGNAL \RegFile[9][0]~q\ : std_logic;
SIGNAL \RegFile[10][0]~feeder_combout\ : std_logic;
SIGNAL \RegFile[10][0]~q\ : std_logic;
SIGNAL \RegFile[8][0]~feeder_combout\ : std_logic;
SIGNAL \RegFile[8][0]~q\ : std_logic;
SIGNAL \Mux90~14_combout\ : std_logic;
SIGNAL \RegFile[12][0]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux90~1_combout\ : std_logic;
SIGNAL \RegFile[23][0]~q\ : std_logic;
SIGNAL \RegFile[21][0]~q\ : std_logic;
SIGNAL \RegFile[22][0]~q\ : std_logic;
SIGNAL \RegFile[19][0]~q\ : std_logic;
SIGNAL \RegFile[18][0]~feeder_combout\ : std_logic;
SIGNAL \RegFile[18][0]~DUPLICATE_q\ : std_logic;
SIGNAL \RegFile[17][0]~q\ : std_logic;
SIGNAL \RegFile[16][0]~q\ : std_logic;
SIGNAL \Mux90~18_combout\ : std_logic;
SIGNAL \RegFile[20][0]~q\ : std_logic;
SIGNAL \Mux90~5_combout\ : std_logic;
SIGNAL \Mux90~13_combout\ : std_logic;
SIGNAL \Mux254~0_combout\ : std_logic;
SIGNAL \Add2~1_OTERM735_OTERM837\ : std_logic;
SIGNAL \Add1~2\ : std_logic;
SIGNAL \Add1~5_sumout\ : std_logic;
SIGNAL \Add2~2\ : std_logic;
SIGNAL \Add2~3\ : std_logic;
SIGNAL \Add2~5_sumout\ : std_logic;
SIGNAL \Mux151~0_combout\ : std_logic;
SIGNAL \RegFile[21][3]~q\ : std_logic;
SIGNAL \RegFile[23][3]~q\ : std_logic;
SIGNAL \RegFile[22][3]~feeder_combout\ : std_logic;
SIGNAL \RegFile[22][3]~q\ : std_logic;
SIGNAL \RegFile[17][3]~q\ : std_logic;
SIGNAL \RegFile[18][3]~q\ : std_logic;
SIGNAL \RegFile[19][3]~feeder_combout\ : std_logic;
SIGNAL \RegFile[19][3]~q\ : std_logic;
SIGNAL \RegFile[16][3]~feeder_combout\ : std_logic;
SIGNAL \RegFile[16][3]~q\ : std_logic;
SIGNAL \Mux87~18_combout\ : std_logic;
SIGNAL \RegFile[20][3]~q\ : std_logic;
SIGNAL \Mux87~5_combout\ : std_logic;
SIGNAL \RegFile[3][3]~q\ : std_logic;
SIGNAL \RegFile[2][3]~q\ : std_logic;
SIGNAL \RegFile[4][3]~feeder_combout\ : std_logic;
SIGNAL \RegFile[4][3]~q\ : std_logic;
SIGNAL \RegFile[5][3]~feeder_combout\ : std_logic;
SIGNAL \RegFile[5][3]~q\ : std_logic;
SIGNAL \RegFile[6][3]~q\ : std_logic;
SIGNAL \RegFile[7][3]~q\ : std_logic;
SIGNAL \Mux87~0_combout\ : std_logic;
SIGNAL \RegFile[1][3]~feeder_combout\ : std_logic;
SIGNAL \RegFile[1][3]~q\ : std_logic;
SIGNAL \Mux87~26_combout\ : std_logic;
SIGNAL \RegFile[15][3]~q\ : std_logic;
SIGNAL \RegFile[14][3]~feeder_combout\ : std_logic;
SIGNAL \RegFile[14][3]~q\ : std_logic;
SIGNAL \RegFile[11][3]~q\ : std_logic;
SIGNAL \RegFile[9][3]~q\ : std_logic;
SIGNAL \RegFile[10][3]~q\ : std_logic;
SIGNAL \RegFile[8][3]~q\ : std_logic;
SIGNAL \Mux87~14_combout\ : std_logic;
SIGNAL \RegFile[12][3]~q\ : std_logic;
SIGNAL \Mux87~1_combout\ : std_logic;
SIGNAL \RegFile[29][3]~q\ : std_logic;
SIGNAL \RegFile[31][3]~q\ : std_logic;
SIGNAL \RegFile[30][3]~q\ : std_logic;
SIGNAL \RegFile[25][3]~q\ : std_logic;
SIGNAL \RegFile[26][3]~q\ : std_logic;
SIGNAL \RegFile[27][3]~q\ : std_logic;
SIGNAL \RegFile[24][3]~feeder_combout\ : std_logic;
SIGNAL \RegFile[24][3]~q\ : std_logic;
SIGNAL \Mux87~22_combout\ : std_logic;
SIGNAL \RegFile[28][3]~feeder_combout\ : std_logic;
SIGNAL \RegFile[28][3]~q\ : std_logic;
SIGNAL \Mux87~9_combout\ : std_logic;
SIGNAL \Mux87~13_combout\ : std_logic;
SIGNAL \Mux251~0_combout\ : std_logic;
SIGNAL \RegFile[13][2]~q\ : std_logic;
SIGNAL \RegFile[14][2]~DUPLICATE_q\ : std_logic;
SIGNAL \RegFile[15][2]~q\ : std_logic;
SIGNAL \RegFile[11][2]~feeder_combout\ : std_logic;
SIGNAL \RegFile[11][2]~q\ : std_logic;
SIGNAL \RegFile[10][2]~feeder_combout\ : std_logic;
SIGNAL \RegFile[10][2]~q\ : std_logic;
SIGNAL \RegFile[9][2]~feeder_combout\ : std_logic;
SIGNAL \RegFile[9][2]~q\ : std_logic;
SIGNAL \RegFile[8][2]~feeder_combout\ : std_logic;
SIGNAL \RegFile[8][2]~q\ : std_logic;
SIGNAL \Mux88~14_combout\ : std_logic;
SIGNAL \RegFile[12][2]~q\ : std_logic;
SIGNAL \Mux88~1_combout\ : std_logic;
SIGNAL \RegFile[31][2]~q\ : std_logic;
SIGNAL \RegFile[29][2]~q\ : std_logic;
SIGNAL \RegFile[30][2]~q\ : std_logic;
SIGNAL \RegFile[27][2]~q\ : std_logic;
SIGNAL \RegFile[25][2]~q\ : std_logic;
SIGNAL \RegFile[26][2]~q\ : std_logic;
SIGNAL \RegFile[24][2]~feeder_combout\ : std_logic;
SIGNAL \RegFile[24][2]~q\ : std_logic;
SIGNAL \Mux88~22_combout\ : std_logic;
SIGNAL \RegFile[28][2]~feeder_combout\ : std_logic;
SIGNAL \RegFile[28][2]~q\ : std_logic;
SIGNAL \Mux88~9_combout\ : std_logic;
SIGNAL \RegFile[21][2]~q\ : std_logic;
SIGNAL \RegFile[23][2]~q\ : std_logic;
SIGNAL \RegFile[22][2]~q\ : std_logic;
SIGNAL \RegFile[17][2]~feeder_combout\ : std_logic;
SIGNAL \RegFile[17][2]~q\ : std_logic;
SIGNAL \RegFile[18][2]~feeder_combout\ : std_logic;
SIGNAL \RegFile[18][2]~q\ : std_logic;
SIGNAL \RegFile[19][2]~feeder_combout\ : std_logic;
SIGNAL \RegFile[19][2]~q\ : std_logic;
SIGNAL \RegFile[16][2]~q\ : std_logic;
SIGNAL \Mux88~18_combout\ : std_logic;
SIGNAL \RegFile[20][2]~q\ : std_logic;
SIGNAL \Mux88~5_combout\ : std_logic;
SIGNAL \RegFile[6][2]~q\ : std_logic;
SIGNAL \RegFile[4][2]~q\ : std_logic;
SIGNAL \RegFile[5][2]~feeder_combout\ : std_logic;
SIGNAL \RegFile[5][2]~q\ : std_logic;
SIGNAL \RegFile[7][2]~q\ : std_logic;
SIGNAL \Mux88~0_combout\ : std_logic;
SIGNAL \RegFile[3][2]~q\ : std_logic;
SIGNAL \RegFile[1][2]~feeder_combout\ : std_logic;
SIGNAL \RegFile[1][2]~q\ : std_logic;
SIGNAL \Mux88~26_combout\ : std_logic;
SIGNAL \Mux88~13_combout\ : std_logic;
SIGNAL \Mux252~0_combout\ : std_logic;
SIGNAL \ShiftLeft0~3_combout\ : std_logic;
SIGNAL \ShiftLeft0~3_OTERM223\ : std_logic;
SIGNAL \R.aluOp.ALUOpXor~DUPLICATE_q\ : std_logic;
SIGNAL \Mux23~0_combout\ : std_logic;
SIGNAL \Mux23~1_combout\ : std_logic;
SIGNAL \R.aluOp.ALUOpXor~q\ : std_logic;
SIGNAL \R.aluOp.ALUOpXor_OTERM355\ : std_logic;
SIGNAL \R.aluOp.ALUOpOr~q\ : std_logic;
SIGNAL \Mux22~0_combout\ : std_logic;
SIGNAL \Mux22~1_combout\ : std_logic;
SIGNAL \R.aluOp.ALUOpOr_OTERM353\ : std_logic;
SIGNAL \R.aluOp.ALUOpAnd~q\ : std_logic;
SIGNAL \R.aluOp.ALUOpAnd~DUPLICATE_q\ : std_logic;
SIGNAL \Mux21~1_combout\ : std_logic;
SIGNAL \Mux21~2_combout\ : std_logic;
SIGNAL \R.aluOp.ALUOpAnd_OTERM357\ : std_logic;
SIGNAL \Selector29~0_RTM0409_combout\ : std_logic;
SIGNAL \Selector29~0_OTERM407\ : std_logic;
SIGNAL \Selector29~1_combout\ : std_logic;
SIGNAL \Mux149~0_combout\ : std_logic;
SIGNAL \Mux123~2_combout\ : std_logic;
SIGNAL \Mux141~0_combout\ : std_logic;
SIGNAL \Mux144~0_combout\ : std_logic;
SIGNAL \Mux130~0_combout\ : std_logic;
SIGNAL \Add2~33_OTERM719_OTERM825\ : std_logic;
SIGNAL \Mux146~0_combout\ : std_logic;
SIGNAL \Mux147~0_combout\ : std_logic;
SIGNAL \Selector17~0_combout\ : std_logic;
SIGNAL \Selector17~0_OTERM391\ : std_logic;
SIGNAL \Mux125~0_combout\ : std_logic;
SIGNAL \Add0~106\ : std_logic;
SIGNAL \Add0~109_sumout\ : std_logic;
SIGNAL \RegFile[13][27]~q\ : std_logic;
SIGNAL \RegFile[15][27]~feeder_combout\ : std_logic;
SIGNAL \RegFile[15][27]~q\ : std_logic;
SIGNAL \RegFile[14][27]~feeder_combout\ : std_logic;
SIGNAL \RegFile[14][27]~q\ : std_logic;
SIGNAL \RegFile[9][27]~q\ : std_logic;
SIGNAL \RegFile[11][27]~q\ : std_logic;
SIGNAL \RegFile[10][27]~q\ : std_logic;
SIGNAL \RegFile[8][27]~q\ : std_logic;
SIGNAL \Mux63~14_combout\ : std_logic;
SIGNAL \RegFile[12][27]~q\ : std_logic;
SIGNAL \Mux63~1_combout\ : std_logic;
SIGNAL \RegFile[23][27]~q\ : std_logic;
SIGNAL \RegFile[22][27]~feeder_combout\ : std_logic;
SIGNAL \RegFile[22][27]~q\ : std_logic;
SIGNAL \RegFile[21][27]~feeder_combout\ : std_logic;
SIGNAL \RegFile[21][27]~q\ : std_logic;
SIGNAL \RegFile[17][27]~q\ : std_logic;
SIGNAL \RegFile[18][27]~feeder_combout\ : std_logic;
SIGNAL \RegFile[18][27]~q\ : std_logic;
SIGNAL \RegFile[19][27]~feeder_combout\ : std_logic;
SIGNAL \RegFile[19][27]~q\ : std_logic;
SIGNAL \RegFile[16][27]~feeder_combout\ : std_logic;
SIGNAL \RegFile[16][27]~q\ : std_logic;
SIGNAL \Mux63~18_combout\ : std_logic;
SIGNAL \RegFile[20][27]~q\ : std_logic;
SIGNAL \Mux63~5_combout\ : std_logic;
SIGNAL \RegFile[4][27]~q\ : std_logic;
SIGNAL \RegFile[6][27]~q\ : std_logic;
SIGNAL \RegFile[5][27]~feeder_combout\ : std_logic;
SIGNAL \RegFile[5][27]~q\ : std_logic;
SIGNAL \RegFile[7][27]~q\ : std_logic;
SIGNAL \Mux63~0_combout\ : std_logic;
SIGNAL \RegFile[3][27]~feeder_combout\ : std_logic;
SIGNAL \RegFile[3][27]~q\ : std_logic;
SIGNAL \RegFile[2][27]~q\ : std_logic;
SIGNAL \RegFile[1][27]~feeder_combout\ : std_logic;
SIGNAL \RegFile[1][27]~q\ : std_logic;
SIGNAL \Mux63~26_combout\ : std_logic;
SIGNAL \RegFile[31][27]~q\ : std_logic;
SIGNAL \RegFile[30][27]~feeder_combout\ : std_logic;
SIGNAL \RegFile[30][27]~q\ : std_logic;
SIGNAL \RegFile[27][27]~q\ : std_logic;
SIGNAL \RegFile[25][27]~q\ : std_logic;
SIGNAL \RegFile[26][27]~feeder_combout\ : std_logic;
SIGNAL \RegFile[26][27]~DUPLICATE_q\ : std_logic;
SIGNAL \RegFile[24][27]~feeder_combout\ : std_logic;
SIGNAL \RegFile[24][27]~q\ : std_logic;
SIGNAL \Mux63~22_combout\ : std_logic;
SIGNAL \RegFile[28][27]~q\ : std_logic;
SIGNAL \Mux63~9_combout\ : std_logic;
SIGNAL \Mux63~13_combout\ : std_logic;
SIGNAL \Mux227~0_combout\ : std_logic;
SIGNAL \Mux128~0_combout\ : std_logic;
SIGNAL \RegFile[3][26]~q\ : std_logic;
SIGNAL \RegFile[2][26]~q\ : std_logic;
SIGNAL \RegFile[7][26]~DUPLICATE_q\ : std_logic;
SIGNAL \RegFile[6][26]~q\ : std_logic;
SIGNAL \RegFile[5][26]~feeder_combout\ : std_logic;
SIGNAL \RegFile[5][26]~q\ : std_logic;
SIGNAL \RegFile[4][26]~feeder_combout\ : std_logic;
SIGNAL \RegFile[4][26]~q\ : std_logic;
SIGNAL \Mux96~0_combout\ : std_logic;
SIGNAL \RegFile[1][26]~feeder_combout\ : std_logic;
SIGNAL \RegFile[1][26]~q\ : std_logic;
SIGNAL \Mux96~26_combout\ : std_logic;
SIGNAL \RegFile[23][26]~q\ : std_logic;
SIGNAL \RegFile[22][26]~q\ : std_logic;
SIGNAL \RegFile[17][26]~q\ : std_logic;
SIGNAL \RegFile[18][26]~feeder_combout\ : std_logic;
SIGNAL \RegFile[18][26]~q\ : std_logic;
SIGNAL \RegFile[19][26]~q\ : std_logic;
SIGNAL \RegFile[16][26]~feeder_combout\ : std_logic;
SIGNAL \RegFile[16][26]~q\ : std_logic;
SIGNAL \Mux96~18_combout\ : std_logic;
SIGNAL \RegFile[20][26]~q\ : std_logic;
SIGNAL \Mux96~5_combout\ : std_logic;
SIGNAL \RegFile[29][26]~q\ : std_logic;
SIGNAL \RegFile[30][26]~feeder_combout\ : std_logic;
SIGNAL \RegFile[30][26]~q\ : std_logic;
SIGNAL \RegFile[31][26]~q\ : std_logic;
SIGNAL \RegFile[25][26]~q\ : std_logic;
SIGNAL \RegFile[26][26]~feeder_combout\ : std_logic;
SIGNAL \RegFile[26][26]~q\ : std_logic;
SIGNAL \RegFile[27][26]~q\ : std_logic;
SIGNAL \RegFile[24][26]~feeder_combout\ : std_logic;
SIGNAL \RegFile[24][26]~q\ : std_logic;
SIGNAL \Mux96~22_combout\ : std_logic;
SIGNAL \RegFile[28][26]~q\ : std_logic;
SIGNAL \Mux96~9_combout\ : std_logic;
SIGNAL \RegFile[15][26]~q\ : std_logic;
SIGNAL \RegFile[14][26]~feeder_combout\ : std_logic;
SIGNAL \RegFile[14][26]~q\ : std_logic;
SIGNAL \RegFile[13][26]~q\ : std_logic;
SIGNAL \RegFile[11][26]~q\ : std_logic;
SIGNAL \RegFile[9][26]~q\ : std_logic;
SIGNAL \RegFile[10][26]~q\ : std_logic;
SIGNAL \RegFile[8][26]~q\ : std_logic;
SIGNAL \Mux96~14_combout\ : std_logic;
SIGNAL \RegFile[12][26]~feeder_combout\ : std_logic;
SIGNAL \RegFile[12][26]~q\ : std_logic;
SIGNAL \Mux96~1_combout\ : std_logic;
SIGNAL \Mux96~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[26]~25_combout\ : std_logic;
SIGNAL \Add0~90\ : std_logic;
SIGNAL \Add0~93_sumout\ : std_logic;
SIGNAL \ShiftRight1~55_combout\ : std_logic;
SIGNAL \Add0~110\ : std_logic;
SIGNAL \Add0~113_sumout\ : std_logic;
SIGNAL \Mux124~1_combout\ : std_logic;
SIGNAL \RegFile[29][30]~q\ : std_logic;
SIGNAL \RegFile[30][30]~feeder_combout\ : std_logic;
SIGNAL \RegFile[30][30]~q\ : std_logic;
SIGNAL \RegFile[31][30]~q\ : std_logic;
SIGNAL \RegFile[27][30]~feeder_combout\ : std_logic;
SIGNAL \RegFile[27][30]~q\ : std_logic;
SIGNAL \RegFile[26][30]~feeder_combout\ : std_logic;
SIGNAL \RegFile[26][30]~q\ : std_logic;
SIGNAL \RegFile[25][30]~q\ : std_logic;
SIGNAL \RegFile[24][30]~q\ : std_logic;
SIGNAL \Mux92~22_combout\ : std_logic;
SIGNAL \RegFile[28][30]~feeder_combout\ : std_logic;
SIGNAL \RegFile[28][30]~q\ : std_logic;
SIGNAL \Mux92~9_combout\ : std_logic;
SIGNAL \RegFile[21][30]~q\ : std_logic;
SIGNAL \RegFile[22][30]~feeder_combout\ : std_logic;
SIGNAL \RegFile[22][30]~q\ : std_logic;
SIGNAL \RegFile[17][30]~q\ : std_logic;
SIGNAL \RegFile[18][30]~feeder_combout\ : std_logic;
SIGNAL \RegFile[18][30]~q\ : std_logic;
SIGNAL \RegFile[19][30]~q\ : std_logic;
SIGNAL \RegFile[16][30]~feeder_combout\ : std_logic;
SIGNAL \RegFile[16][30]~q\ : std_logic;
SIGNAL \Mux92~18_combout\ : std_logic;
SIGNAL \RegFile[20][30]~feeder_combout\ : std_logic;
SIGNAL \RegFile[20][30]~q\ : std_logic;
SIGNAL \Mux92~5_combout\ : std_logic;
SIGNAL \RegFile[3][30]~q\ : std_logic;
SIGNAL \RegFile[2][30]~q\ : std_logic;
SIGNAL \RegFile[6][30]~q\ : std_logic;
SIGNAL \RegFile[4][30]~q\ : std_logic;
SIGNAL \RegFile[7][30]~q\ : std_logic;
SIGNAL \RegFile[5][30]~q\ : std_logic;
SIGNAL \Mux92~0_combout\ : std_logic;
SIGNAL \RegFile[1][30]~feeder_combout\ : std_logic;
SIGNAL \RegFile[1][30]~q\ : std_logic;
SIGNAL \Mux92~26_combout\ : std_logic;
SIGNAL \RegFile[13][30]~q\ : std_logic;
SIGNAL \RegFile[15][30]~q\ : std_logic;
SIGNAL \RegFile[14][30]~q\ : std_logic;
SIGNAL \RegFile[11][30]~q\ : std_logic;
SIGNAL \RegFile[9][30]~q\ : std_logic;
SIGNAL \RegFile[10][30]~feeder_combout\ : std_logic;
SIGNAL \RegFile[10][30]~q\ : std_logic;
SIGNAL \RegFile[8][30]~feeder_combout\ : std_logic;
SIGNAL \RegFile[8][30]~q\ : std_logic;
SIGNAL \Mux92~14_combout\ : std_logic;
SIGNAL \RegFile[12][30]~q\ : std_logic;
SIGNAL \Mux92~1_combout\ : std_logic;
SIGNAL \Mux92~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[30]~30_combout\ : std_logic;
SIGNAL \Add1~118\ : std_logic;
SIGNAL \Add1~121_sumout\ : std_logic;
SIGNAL \Mux129~0_combout\ : std_logic;
SIGNAL \RegFile[2][25]~q\ : std_logic;
SIGNAL \RegFile[3][25]~q\ : std_logic;
SIGNAL \RegFile[6][25]~q\ : std_logic;
SIGNAL \RegFile[7][25]~q\ : std_logic;
SIGNAL \RegFile[4][25]~feeder_combout\ : std_logic;
SIGNAL \RegFile[4][25]~q\ : std_logic;
SIGNAL \RegFile[5][25]~feeder_combout\ : std_logic;
SIGNAL \RegFile[5][25]~q\ : std_logic;
SIGNAL \Mux97~0_combout\ : std_logic;
SIGNAL \RegFile[1][25]~q\ : std_logic;
SIGNAL \Mux97~26_combout\ : std_logic;
SIGNAL \RegFile[30][25]~feeder_combout\ : std_logic;
SIGNAL \RegFile[30][25]~q\ : std_logic;
SIGNAL \RegFile[29][25]~q\ : std_logic;
SIGNAL \RegFile[25][25]~q\ : std_logic;
SIGNAL \RegFile[26][25]~q\ : std_logic;
SIGNAL \RegFile[27][25]~q\ : std_logic;
SIGNAL \RegFile[24][25]~feeder_combout\ : std_logic;
SIGNAL \RegFile[24][25]~q\ : std_logic;
SIGNAL \Mux97~22_combout\ : std_logic;
SIGNAL \RegFile[28][25]~feeder_combout\ : std_logic;
SIGNAL \RegFile[28][25]~q\ : std_logic;
SIGNAL \Mux97~9_combout\ : std_logic;
SIGNAL \RegFile[15][25]~q\ : std_logic;
SIGNAL \RegFile[13][25]~q\ : std_logic;
SIGNAL \RegFile[14][25]~feeder_combout\ : std_logic;
SIGNAL \RegFile[14][25]~q\ : std_logic;
SIGNAL \RegFile[11][25]~q\ : std_logic;
SIGNAL \RegFile[9][25]~q\ : std_logic;
SIGNAL \RegFile[10][25]~q\ : std_logic;
SIGNAL \RegFile[8][25]~q\ : std_logic;
SIGNAL \Mux97~14_combout\ : std_logic;
SIGNAL \RegFile[12][25]~feeder_combout\ : std_logic;
SIGNAL \RegFile[12][25]~q\ : std_logic;
SIGNAL \Mux97~1_combout\ : std_logic;
SIGNAL \RegFile[21][25]~q\ : std_logic;
SIGNAL \RegFile[22][25]~q\ : std_logic;
SIGNAL \RegFile[23][25]~q\ : std_logic;
SIGNAL \RegFile[17][25]~q\ : std_logic;
SIGNAL \RegFile[19][25]~q\ : std_logic;
SIGNAL \RegFile[18][25]~feeder_combout\ : std_logic;
SIGNAL \RegFile[18][25]~q\ : std_logic;
SIGNAL \RegFile[16][25]~feeder_combout\ : std_logic;
SIGNAL \RegFile[16][25]~q\ : std_logic;
SIGNAL \Mux97~18_combout\ : std_logic;
SIGNAL \RegFile[20][25]~feeder_combout\ : std_logic;
SIGNAL \RegFile[20][25]~q\ : std_logic;
SIGNAL \Mux97~5_combout\ : std_logic;
SIGNAL \Mux97~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[25]~22_combout\ : std_logic;
SIGNAL \R.aluData2[25]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux134~0_combout\ : std_logic;
SIGNAL \Add0~73_sumout\ : std_logic;
SIGNAL \R.regWriteData[20]~feeder_combout\ : std_logic;
SIGNAL \ShiftRight0~7_RTM0235_combout\ : std_logic;
SIGNAL \ShiftRight0~7_OTERM233DUPLICATE_q\ : std_logic;
SIGNAL \ShiftLeft0~4_combout\ : std_logic;
SIGNAL \ShiftLeft0~4_OTERM237\ : std_logic;
SIGNAL \Selector12~3_combout\ : std_logic;
SIGNAL \Selector12~4_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[20]~3_combout\ : std_logic;
SIGNAL \Mux137~0_combout\ : std_logic;
SIGNAL \Mux139~0_combout\ : std_logic;
SIGNAL \Add0~46\ : std_logic;
SIGNAL \Add0~50\ : std_logic;
SIGNAL \Add0~53_sumout\ : std_logic;
SIGNAL \R.regWriteData[15]~feeder_combout\ : std_logic;
SIGNAL \RegFile[29][15]~q\ : std_logic;
SIGNAL \RegFile[30][15]~q\ : std_logic;
SIGNAL \RegFile[27][15]~q\ : std_logic;
SIGNAL \RegFile[26][15]~q\ : std_logic;
SIGNAL \RegFile[25][15]~q\ : std_logic;
SIGNAL \RegFile[24][15]~q\ : std_logic;
SIGNAL \Mux75~22_combout\ : std_logic;
SIGNAL \RegFile[28][15]~q\ : std_logic;
SIGNAL \Mux75~9_combout\ : std_logic;
SIGNAL \RegFile[15][15]~q\ : std_logic;
SIGNAL \RegFile[14][15]~q\ : std_logic;
SIGNAL \RegFile[13][15]~q\ : std_logic;
SIGNAL \RegFile[11][15]~q\ : std_logic;
SIGNAL \RegFile[10][15]~q\ : std_logic;
SIGNAL \RegFile[9][15]~q\ : std_logic;
SIGNAL \RegFile[8][15]~q\ : std_logic;
SIGNAL \Mux75~14_combout\ : std_logic;
SIGNAL \RegFile[12][15]~feeder_combout\ : std_logic;
SIGNAL \RegFile[12][15]~q\ : std_logic;
SIGNAL \Mux75~1_combout\ : std_logic;
SIGNAL \RegFile[3][15]~q\ : std_logic;
SIGNAL \RegFile[2][15]~q\ : std_logic;
SIGNAL \RegFile[4][15]~feeder_combout\ : std_logic;
SIGNAL \RegFile[4][15]~q\ : std_logic;
SIGNAL \RegFile[6][15]~q\ : std_logic;
SIGNAL \RegFile[5][15]~q\ : std_logic;
SIGNAL \RegFile[7][15]~q\ : std_logic;
SIGNAL \Mux75~0_combout\ : std_logic;
SIGNAL \RegFile[1][15]~q\ : std_logic;
SIGNAL \Mux75~26_combout\ : std_logic;
SIGNAL \RegFile[23][15]~q\ : std_logic;
SIGNAL \RegFile[22][15]~feeder_combout\ : std_logic;
SIGNAL \RegFile[22][15]~q\ : std_logic;
SIGNAL \RegFile[21][15]~q\ : std_logic;
SIGNAL \RegFile[17][15]~feeder_combout\ : std_logic;
SIGNAL \RegFile[17][15]~q\ : std_logic;
SIGNAL \RegFile[18][15]~feeder_combout\ : std_logic;
SIGNAL \RegFile[18][15]~q\ : std_logic;
SIGNAL \RegFile[19][15]~q\ : std_logic;
SIGNAL \RegFile[16][15]~feeder_combout\ : std_logic;
SIGNAL \RegFile[16][15]~q\ : std_logic;
SIGNAL \Mux75~18_combout\ : std_logic;
SIGNAL \RegFile[20][15]~q\ : std_logic;
SIGNAL \Mux75~5_combout\ : std_logic;
SIGNAL \Mux75~13_combout\ : std_logic;
SIGNAL \Mux239~0_combout\ : std_logic;
SIGNAL \Mux140~0_combout\ : std_logic;
SIGNAL \Add0~49_sumout\ : std_logic;
SIGNAL \R.regWriteData[14]~feeder_combout\ : std_logic;
SIGNAL \Add2~57_OTERM707_OTERM813\ : std_logic;
SIGNAL \Mux142~0_combout\ : std_logic;
SIGNAL \RegFile[31][12]~q\ : std_logic;
SIGNAL \RegFile[29][12]~q\ : std_logic;
SIGNAL \RegFile[30][12]~q\ : std_logic;
SIGNAL \RegFile[25][12]~q\ : std_logic;
SIGNAL \RegFile[26][12]~feeder_combout\ : std_logic;
SIGNAL \RegFile[26][12]~q\ : std_logic;
SIGNAL \RegFile[27][12]~q\ : std_logic;
SIGNAL \RegFile[24][12]~feeder_combout\ : std_logic;
SIGNAL \RegFile[24][12]~q\ : std_logic;
SIGNAL \Mux110~22_combout\ : std_logic;
SIGNAL \RegFile[28][12]~feeder_combout\ : std_logic;
SIGNAL \RegFile[28][12]~q\ : std_logic;
SIGNAL \Mux110~9_combout\ : std_logic;
SIGNAL \RegFile[3][12]~feeder_combout\ : std_logic;
SIGNAL \RegFile[3][12]~q\ : std_logic;
SIGNAL \RegFile[2][12]~q\ : std_logic;
SIGNAL \RegFile[5][12]~q\ : std_logic;
SIGNAL \RegFile[7][12]~q\ : std_logic;
SIGNAL \RegFile[4][12]~q\ : std_logic;
SIGNAL \RegFile[6][12]~q\ : std_logic;
SIGNAL \Mux110~0_combout\ : std_logic;
SIGNAL \RegFile[1][12]~feeder_combout\ : std_logic;
SIGNAL \RegFile[1][12]~q\ : std_logic;
SIGNAL \Mux110~26_combout\ : std_logic;
SIGNAL \RegFile[21][12]~q\ : std_logic;
SIGNAL \RegFile[23][12]~q\ : std_logic;
SIGNAL \RegFile[22][12]~q\ : std_logic;
SIGNAL \RegFile[17][12]~q\ : std_logic;
SIGNAL \RegFile[18][12]~feeder_combout\ : std_logic;
SIGNAL \RegFile[18][12]~q\ : std_logic;
SIGNAL \RegFile[19][12]~q\ : std_logic;
SIGNAL \RegFile[16][12]~q\ : std_logic;
SIGNAL \Mux110~18_combout\ : std_logic;
SIGNAL \RegFile[20][12]~feeder_combout\ : std_logic;
SIGNAL \RegFile[20][12]~q\ : std_logic;
SIGNAL \Mux110~5_combout\ : std_logic;
SIGNAL \RegFile[15][12]~q\ : std_logic;
SIGNAL \RegFile[14][12]~q\ : std_logic;
SIGNAL \RegFile[9][12]~q\ : std_logic;
SIGNAL \RegFile[10][12]~feeder_combout\ : std_logic;
SIGNAL \RegFile[10][12]~q\ : std_logic;
SIGNAL \RegFile[11][12]~q\ : std_logic;
SIGNAL \RegFile[8][12]~q\ : std_logic;
SIGNAL \Mux110~14_combout\ : std_logic;
SIGNAL \RegFile[12][12]~feeder_combout\ : std_logic;
SIGNAL \RegFile[12][12]~q\ : std_logic;
SIGNAL \Mux110~1_combout\ : std_logic;
SIGNAL \Mux110~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[12]~11_combout\ : std_logic;
SIGNAL \Mux143~0_combout\ : std_logic;
SIGNAL \Mux143~1_combout\ : std_logic;
SIGNAL \RegFile[31][11]~q\ : std_logic;
SIGNAL \RegFile[30][11]~q\ : std_logic;
SIGNAL \RegFile[25][11]~q\ : std_logic;
SIGNAL \RegFile[27][11]~feeder_combout\ : std_logic;
SIGNAL \RegFile[27][11]~q\ : std_logic;
SIGNAL \RegFile[26][11]~feeder_combout\ : std_logic;
SIGNAL \RegFile[26][11]~q\ : std_logic;
SIGNAL \RegFile[24][11]~feeder_combout\ : std_logic;
SIGNAL \RegFile[24][11]~q\ : std_logic;
SIGNAL \Mux111~22_combout\ : std_logic;
SIGNAL \RegFile[28][11]~feeder_combout\ : std_logic;
SIGNAL \RegFile[28][11]~q\ : std_logic;
SIGNAL \Mux111~9_combout\ : std_logic;
SIGNAL \RegFile[15][11]~feeder_combout\ : std_logic;
SIGNAL \RegFile[15][11]~q\ : std_logic;
SIGNAL \RegFile[13][11]~q\ : std_logic;
SIGNAL \RegFile[14][11]~feeder_combout\ : std_logic;
SIGNAL \RegFile[14][11]~q\ : std_logic;
SIGNAL \RegFile[9][11]~q\ : std_logic;
SIGNAL \RegFile[11][11]~feeder_combout\ : std_logic;
SIGNAL \RegFile[11][11]~DUPLICATE_q\ : std_logic;
SIGNAL \RegFile[10][11]~feeder_combout\ : std_logic;
SIGNAL \RegFile[10][11]~q\ : std_logic;
SIGNAL \RegFile[8][11]~feeder_combout\ : std_logic;
SIGNAL \RegFile[8][11]~q\ : std_logic;
SIGNAL \Mux111~14_combout\ : std_logic;
SIGNAL \RegFile[12][11]~q\ : std_logic;
SIGNAL \Mux111~1_combout\ : std_logic;
SIGNAL \RegFile[21][11]~q\ : std_logic;
SIGNAL \RegFile[23][11]~q\ : std_logic;
SIGNAL \RegFile[22][11]~feeder_combout\ : std_logic;
SIGNAL \RegFile[22][11]~q\ : std_logic;
SIGNAL \RegFile[19][11]~q\ : std_logic;
SIGNAL \RegFile[17][11]~q\ : std_logic;
SIGNAL \RegFile[18][11]~q\ : std_logic;
SIGNAL \RegFile[16][11]~q\ : std_logic;
SIGNAL \Mux111~18_combout\ : std_logic;
SIGNAL \RegFile[20][11]~feeder_combout\ : std_logic;
SIGNAL \RegFile[20][11]~q\ : std_logic;
SIGNAL \Mux111~5_combout\ : std_logic;
SIGNAL \RegFile[3][11]~q\ : std_logic;
SIGNAL \RegFile[2][11]~q\ : std_logic;
SIGNAL \RegFile[6][11]~q\ : std_logic;
SIGNAL \RegFile[7][11]~q\ : std_logic;
SIGNAL \RegFile[4][11]~feeder_combout\ : std_logic;
SIGNAL \RegFile[4][11]~q\ : std_logic;
SIGNAL \RegFile[5][11]~q\ : std_logic;
SIGNAL \Mux111~0_combout\ : std_logic;
SIGNAL \RegFile[1][11]~feeder_combout\ : std_logic;
SIGNAL \RegFile[1][11]~q\ : std_logic;
SIGNAL \Mux111~26_combout\ : std_logic;
SIGNAL \Mux111~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[11]~8_combout\ : std_logic;
SIGNAL \Add2~41_OTERM715_OTERM819\ : std_logic;
SIGNAL \RegFile[13][10]~feeder_combout\ : std_logic;
SIGNAL \RegFile[13][10]~q\ : std_logic;
SIGNAL \RegFile[14][10]~feeder_combout\ : std_logic;
SIGNAL \RegFile[14][10]~q\ : std_logic;
SIGNAL \RegFile[15][10]~q\ : std_logic;
SIGNAL \RegFile[9][10]~feeder_combout\ : std_logic;
SIGNAL \RegFile[9][10]~q\ : std_logic;
SIGNAL \RegFile[11][10]~q\ : std_logic;
SIGNAL \RegFile[10][10]~feeder_combout\ : std_logic;
SIGNAL \RegFile[10][10]~q\ : std_logic;
SIGNAL \RegFile[8][10]~feeder_combout\ : std_logic;
SIGNAL \RegFile[8][10]~q\ : std_logic;
SIGNAL \Mux80~14_combout\ : std_logic;
SIGNAL \RegFile[12][10]~feeder_combout\ : std_logic;
SIGNAL \RegFile[12][10]~q\ : std_logic;
SIGNAL \Mux80~1_combout\ : std_logic;
SIGNAL \RegFile[31][10]~q\ : std_logic;
SIGNAL \RegFile[30][10]~q\ : std_logic;
SIGNAL \RegFile[29][10]~q\ : std_logic;
SIGNAL \RegFile[27][10]~q\ : std_logic;
SIGNAL \RegFile[26][10]~q\ : std_logic;
SIGNAL \RegFile[25][10]~q\ : std_logic;
SIGNAL \RegFile[24][10]~q\ : std_logic;
SIGNAL \Mux80~22_combout\ : std_logic;
SIGNAL \RegFile[28][10]~q\ : std_logic;
SIGNAL \Mux80~9_combout\ : std_logic;
SIGNAL \RegFile[21][10]~q\ : std_logic;
SIGNAL \RegFile[23][10]~q\ : std_logic;
SIGNAL \RegFile[22][10]~q\ : std_logic;
SIGNAL \RegFile[17][10]~q\ : std_logic;
SIGNAL \RegFile[18][10]~q\ : std_logic;
SIGNAL \RegFile[19][10]~feeder_combout\ : std_logic;
SIGNAL \RegFile[19][10]~q\ : std_logic;
SIGNAL \RegFile[16][10]~feeder_combout\ : std_logic;
SIGNAL \RegFile[16][10]~q\ : std_logic;
SIGNAL \Mux80~18_combout\ : std_logic;
SIGNAL \RegFile[20][10]~q\ : std_logic;
SIGNAL \Mux80~5_combout\ : std_logic;
SIGNAL \RegFile[3][10]~q\ : std_logic;
SIGNAL \RegFile[6][10]~q\ : std_logic;
SIGNAL \RegFile[5][10]~feeder_combout\ : std_logic;
SIGNAL \RegFile[5][10]~q\ : std_logic;
SIGNAL \RegFile[7][10]~q\ : std_logic;
SIGNAL \RegFile[4][10]~q\ : std_logic;
SIGNAL \Mux80~0_combout\ : std_logic;
SIGNAL \RegFile[1][10]~feeder_combout\ : std_logic;
SIGNAL \RegFile[1][10]~q\ : std_logic;
SIGNAL \Mux80~26_combout\ : std_logic;
SIGNAL \Mux80~13_combout\ : std_logic;
SIGNAL \Mux244~0_combout\ : std_logic;
SIGNAL \Add2~41_OTERM715_OTERM817feeder_combout\ : std_logic;
SIGNAL \Add2~41_OTERM715_OTERM817\ : std_logic;
SIGNAL \Mux145~0_combout\ : std_logic;
SIGNAL \Add0~26\ : std_logic;
SIGNAL \Add0~29_sumout\ : std_logic;
SIGNAL \R.regWriteData[9]~feeder_combout\ : std_logic;
SIGNAL \RegFile[31][9]~feeder_combout\ : std_logic;
SIGNAL \RegFile[31][9]~q\ : std_logic;
SIGNAL \RegFile[30][9]~feeder_combout\ : std_logic;
SIGNAL \RegFile[30][9]~q\ : std_logic;
SIGNAL \RegFile[29][9]~feeder_combout\ : std_logic;
SIGNAL \RegFile[29][9]~q\ : std_logic;
SIGNAL \RegFile[25][9]~q\ : std_logic;
SIGNAL \RegFile[26][9]~feeder_combout\ : std_logic;
SIGNAL \RegFile[26][9]~q\ : std_logic;
SIGNAL \RegFile[27][9]~q\ : std_logic;
SIGNAL \RegFile[24][9]~q\ : std_logic;
SIGNAL \Mux81~22_combout\ : std_logic;
SIGNAL \RegFile[28][9]~q\ : std_logic;
SIGNAL \Mux81~9_combout\ : std_logic;
SIGNAL \RegFile[14][9]~q\ : std_logic;
SIGNAL \RegFile[15][9]~q\ : std_logic;
SIGNAL \RegFile[9][9]~q\ : std_logic;
SIGNAL \RegFile[10][9]~q\ : std_logic;
SIGNAL \RegFile[11][9]~q\ : std_logic;
SIGNAL \RegFile[8][9]~feeder_combout\ : std_logic;
SIGNAL \RegFile[8][9]~q\ : std_logic;
SIGNAL \Mux81~14_combout\ : std_logic;
SIGNAL \RegFile[12][9]~feeder_combout\ : std_logic;
SIGNAL \RegFile[12][9]~q\ : std_logic;
SIGNAL \Mux81~1_combout\ : std_logic;
SIGNAL \RegFile[23][9]~q\ : std_logic;
SIGNAL \RegFile[21][9]~q\ : std_logic;
SIGNAL \RegFile[22][9]~feeder_combout\ : std_logic;
SIGNAL \RegFile[22][9]~DUPLICATE_q\ : std_logic;
SIGNAL \RegFile[17][9]~DUPLICATE_q\ : std_logic;
SIGNAL \RegFile[18][9]~feeder_combout\ : std_logic;
SIGNAL \RegFile[18][9]~q\ : std_logic;
SIGNAL \RegFile[19][9]~q\ : std_logic;
SIGNAL \RegFile[16][9]~feeder_combout\ : std_logic;
SIGNAL \RegFile[16][9]~q\ : std_logic;
SIGNAL \Mux81~18_combout\ : std_logic;
SIGNAL \RegFile[20][9]~q\ : std_logic;
SIGNAL \Mux81~5_combout\ : std_logic;
SIGNAL \RegFile[3][9]~q\ : std_logic;
SIGNAL \RegFile[2][9]~q\ : std_logic;
SIGNAL \RegFile[6][9]~q\ : std_logic;
SIGNAL \RegFile[5][9]~q\ : std_logic;
SIGNAL \RegFile[4][9]~q\ : std_logic;
SIGNAL \RegFile[7][9]~q\ : std_logic;
SIGNAL \Mux81~0_combout\ : std_logic;
SIGNAL \RegFile[1][9]~q\ : std_logic;
SIGNAL \Mux81~26_combout\ : std_logic;
SIGNAL \Mux81~13_combout\ : std_logic;
SIGNAL \Mux245~0_combout\ : std_logic;
SIGNAL \Add2~33_OTERM719_OTERM821\ : std_logic;
SIGNAL \RegFile[29][7]~q\ : std_logic;
SIGNAL \RegFile[31][7]~q\ : std_logic;
SIGNAL \RegFile[30][7]~feeder_combout\ : std_logic;
SIGNAL \RegFile[30][7]~DUPLICATE_q\ : std_logic;
SIGNAL \RegFile[25][7]~q\ : std_logic;
SIGNAL \RegFile[26][7]~q\ : std_logic;
SIGNAL \RegFile[27][7]~q\ : std_logic;
SIGNAL \RegFile[24][7]~feeder_combout\ : std_logic;
SIGNAL \RegFile[24][7]~q\ : std_logic;
SIGNAL \Mux83~22_combout\ : std_logic;
SIGNAL \RegFile[28][7]~feeder_combout\ : std_logic;
SIGNAL \RegFile[28][7]~q\ : std_logic;
SIGNAL \Mux83~9_combout\ : std_logic;
SIGNAL \RegFile[3][7]~q\ : std_logic;
SIGNAL \RegFile[2][7]~DUPLICATE_q\ : std_logic;
SIGNAL \RegFile[4][7]~feeder_combout\ : std_logic;
SIGNAL \RegFile[4][7]~q\ : std_logic;
SIGNAL \RegFile[6][7]~feeder_combout\ : std_logic;
SIGNAL \RegFile[6][7]~q\ : std_logic;
SIGNAL \RegFile[5][7]~q\ : std_logic;
SIGNAL \RegFile[7][7]~q\ : std_logic;
SIGNAL \Mux83~0_combout\ : std_logic;
SIGNAL \RegFile[1][7]~feeder_combout\ : std_logic;
SIGNAL \RegFile[1][7]~q\ : std_logic;
SIGNAL \Mux83~26_combout\ : std_logic;
SIGNAL \RegFile[21][7]~q\ : std_logic;
SIGNAL \RegFile[22][7]~feeder_combout\ : std_logic;
SIGNAL \RegFile[22][7]~q\ : std_logic;
SIGNAL \RegFile[23][7]~q\ : std_logic;
SIGNAL \RegFile[17][7]~q\ : std_logic;
SIGNAL \RegFile[18][7]~q\ : std_logic;
SIGNAL \RegFile[19][7]~q\ : std_logic;
SIGNAL \RegFile[16][7]~feeder_combout\ : std_logic;
SIGNAL \RegFile[16][7]~q\ : std_logic;
SIGNAL \Mux83~18_combout\ : std_logic;
SIGNAL \RegFile[20][7]~q\ : std_logic;
SIGNAL \Mux83~5_combout\ : std_logic;
SIGNAL \RegFile[15][7]~q\ : std_logic;
SIGNAL \RegFile[14][7]~q\ : std_logic;
SIGNAL \RegFile[13][7]~q\ : std_logic;
SIGNAL \RegFile[11][7]~q\ : std_logic;
SIGNAL \RegFile[9][7]~feeder_combout\ : std_logic;
SIGNAL \RegFile[9][7]~q\ : std_logic;
SIGNAL \RegFile[10][7]~q\ : std_logic;
SIGNAL \RegFile[8][7]~feeder_combout\ : std_logic;
SIGNAL \RegFile[8][7]~q\ : std_logic;
SIGNAL \Mux83~14_combout\ : std_logic;
SIGNAL \RegFile[12][7]~q\ : std_logic;
SIGNAL \Mux83~1_combout\ : std_logic;
SIGNAL \Mux83~13_combout\ : std_logic;
SIGNAL \Mux247~0_combout\ : std_logic;
SIGNAL \Add2~25_OTERM723_OTERM829\ : std_logic;
SIGNAL \Mux148~0_combout\ : std_logic;
SIGNAL \Add0~17_sumout\ : std_logic;
SIGNAL \R.regWriteData[6]~feeder_combout\ : std_logic;
SIGNAL \Selector26~2_RTM0417_combout\ : std_logic;
SIGNAL \Selector26~2_OTERM415\ : std_logic;
SIGNAL \ShiftLeft0~2_combout\ : std_logic;
SIGNAL \ShiftLeft0~2_OTERM221\ : std_logic;
SIGNAL \Selector27~0_combout\ : std_logic;
SIGNAL \Selector27~0_OTERM385\ : std_logic;
SIGNAL \RegFile[21][4]~q\ : std_logic;
SIGNAL \RegFile[22][4]~q\ : std_logic;
SIGNAL \RegFile[17][4]~q\ : std_logic;
SIGNAL \RegFile[18][4]~feeder_combout\ : std_logic;
SIGNAL \RegFile[18][4]~q\ : std_logic;
SIGNAL \RegFile[19][4]~q\ : std_logic;
SIGNAL \RegFile[16][4]~q\ : std_logic;
SIGNAL \Mux86~18_combout\ : std_logic;
SIGNAL \RegFile[20][4]~feeder_combout\ : std_logic;
SIGNAL \RegFile[20][4]~q\ : std_logic;
SIGNAL \Mux86~5_combout\ : std_logic;
SIGNAL \RegFile[31][4]~q\ : std_logic;
SIGNAL \RegFile[29][4]~q\ : std_logic;
SIGNAL \RegFile[30][4]~feeder_combout\ : std_logic;
SIGNAL \RegFile[30][4]~q\ : std_logic;
SIGNAL \RegFile[25][4]~q\ : std_logic;
SIGNAL \RegFile[27][4]~q\ : std_logic;
SIGNAL \RegFile[26][4]~feeder_combout\ : std_logic;
SIGNAL \RegFile[26][4]~q\ : std_logic;
SIGNAL \RegFile[24][4]~feeder_combout\ : std_logic;
SIGNAL \RegFile[24][4]~q\ : std_logic;
SIGNAL \Mux86~22_combout\ : std_logic;
SIGNAL \RegFile[28][4]~feeder_combout\ : std_logic;
SIGNAL \RegFile[28][4]~q\ : std_logic;
SIGNAL \Mux86~9_combout\ : std_logic;
SIGNAL \RegFile[2][4]~q\ : std_logic;
SIGNAL \RegFile[3][4]~feeder_combout\ : std_logic;
SIGNAL \RegFile[3][4]~q\ : std_logic;
SIGNAL \RegFile[5][4]~q\ : std_logic;
SIGNAL \RegFile[6][4]~feeder_combout\ : std_logic;
SIGNAL \RegFile[6][4]~q\ : std_logic;
SIGNAL \RegFile[4][4]~feeder_combout\ : std_logic;
SIGNAL \RegFile[4][4]~q\ : std_logic;
SIGNAL \RegFile[7][4]~q\ : std_logic;
SIGNAL \Mux86~0_combout\ : std_logic;
SIGNAL \RegFile[1][4]~feeder_combout\ : std_logic;
SIGNAL \RegFile[1][4]~q\ : std_logic;
SIGNAL \Mux86~26_combout\ : std_logic;
SIGNAL \RegFile[13][4]~q\ : std_logic;
SIGNAL \RegFile[14][4]~feeder_combout\ : std_logic;
SIGNAL \RegFile[14][4]~q\ : std_logic;
SIGNAL \RegFile[15][4]~q\ : std_logic;
SIGNAL \RegFile[11][4]~q\ : std_logic;
SIGNAL \RegFile[10][4]~feeder_combout\ : std_logic;
SIGNAL \RegFile[10][4]~q\ : std_logic;
SIGNAL \RegFile[9][4]~q\ : std_logic;
SIGNAL \RegFile[8][4]~feeder_combout\ : std_logic;
SIGNAL \RegFile[8][4]~q\ : std_logic;
SIGNAL \Mux86~14_combout\ : std_logic;
SIGNAL \RegFile[12][4]~q\ : std_logic;
SIGNAL \Mux86~1_combout\ : std_logic;
SIGNAL \Mux86~13_combout\ : std_logic;
SIGNAL \Mux250~0_combout\ : std_logic;
SIGNAL \Add0~2\ : std_logic;
SIGNAL \Add0~6\ : std_logic;
SIGNAL \Add0~10\ : std_logic;
SIGNAL \Add0~13_sumout\ : std_logic;
SIGNAL \R.regWriteData[5]~feeder_combout\ : std_logic;
SIGNAL \avm_d_readdata[29]~input_o\ : std_logic;
SIGNAL \ShiftLeft0~7_combout\ : std_logic;
SIGNAL \ShiftLeft0~7_OTERM205\ : std_logic;
SIGNAL \Mux149~1_combout\ : std_logic;
SIGNAL \RegFile[15][5]~q\ : std_logic;
SIGNAL \RegFile[13][5]~q\ : std_logic;
SIGNAL \RegFile[14][5]~feeder_combout\ : std_logic;
SIGNAL \RegFile[14][5]~q\ : std_logic;
SIGNAL \RegFile[11][5]~q\ : std_logic;
SIGNAL \RegFile[10][5]~feeder_combout\ : std_logic;
SIGNAL \RegFile[10][5]~q\ : std_logic;
SIGNAL \RegFile[9][5]~q\ : std_logic;
SIGNAL \RegFile[8][5]~q\ : std_logic;
SIGNAL \Mux117~14_combout\ : std_logic;
SIGNAL \RegFile[12][5]~q\ : std_logic;
SIGNAL \Mux117~1_combout\ : std_logic;
SIGNAL \RegFile[3][5]~q\ : std_logic;
SIGNAL \RegFile[2][5]~q\ : std_logic;
SIGNAL \RegFile[4][5]~feeder_combout\ : std_logic;
SIGNAL \RegFile[4][5]~q\ : std_logic;
SIGNAL \RegFile[7][5]~q\ : std_logic;
SIGNAL \RegFile[5][5]~q\ : std_logic;
SIGNAL \RegFile[6][5]~q\ : std_logic;
SIGNAL \Mux117~0_combout\ : std_logic;
SIGNAL \RegFile[1][5]~feeder_combout\ : std_logic;
SIGNAL \RegFile[1][5]~q\ : std_logic;
SIGNAL \Mux117~26_combout\ : std_logic;
SIGNAL \RegFile[21][5]~q\ : std_logic;
SIGNAL \RegFile[23][5]~feeder_combout\ : std_logic;
SIGNAL \RegFile[23][5]~q\ : std_logic;
SIGNAL \RegFile[22][5]~feeder_combout\ : std_logic;
SIGNAL \RegFile[22][5]~q\ : std_logic;
SIGNAL \RegFile[19][5]~q\ : std_logic;
SIGNAL \RegFile[18][5]~q\ : std_logic;
SIGNAL \RegFile[17][5]~q\ : std_logic;
SIGNAL \RegFile[16][5]~feeder_combout\ : std_logic;
SIGNAL \RegFile[16][5]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux117~18_combout\ : std_logic;
SIGNAL \RegFile[20][5]~feeder_combout\ : std_logic;
SIGNAL \RegFile[20][5]~q\ : std_logic;
SIGNAL \Mux117~5_combout\ : std_logic;
SIGNAL \RegFile[31][5]~q\ : std_logic;
SIGNAL \RegFile[30][5]~q\ : std_logic;
SIGNAL \RegFile[27][5]~feeder_combout\ : std_logic;
SIGNAL \RegFile[27][5]~q\ : std_logic;
SIGNAL \RegFile[25][5]~feeder_combout\ : std_logic;
SIGNAL \RegFile[25][5]~q\ : std_logic;
SIGNAL \RegFile[26][5]~feeder_combout\ : std_logic;
SIGNAL \RegFile[26][5]~q\ : std_logic;
SIGNAL \RegFile[24][5]~feeder_combout\ : std_logic;
SIGNAL \RegFile[24][5]~q\ : std_logic;
SIGNAL \Mux117~22_combout\ : std_logic;
SIGNAL \RegFile[28][5]~q\ : std_logic;
SIGNAL \Mux117~9_combout\ : std_logic;
SIGNAL \Mux117~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[5]~21_combout\ : std_logic;
SIGNAL \Selector27~2_RTM0413_combout\ : std_logic;
SIGNAL \Selector27~2_OTERM411\ : std_logic;
SIGNAL \ShiftLeft0~6_combout\ : std_logic;
SIGNAL \ShiftLeft0~6_OTERM243\ : std_logic;
SIGNAL \Selector27~3_combout\ : std_logic;
SIGNAL \ShiftRight1~11_combout\ : std_logic;
SIGNAL \ShiftRight1~11_OTERM35\ : std_logic;
SIGNAL \ShiftRight0~8_combout\ : std_logic;
SIGNAL \ShiftRight1~16_combout\ : std_logic;
SIGNAL \ShiftRight1~16_OTERM209\ : std_logic;
SIGNAL \ShiftRight1~17_combout\ : std_logic;
SIGNAL \ShiftRight1~17_OTERM267\ : std_logic;
SIGNAL \RegFile[3][17]~q\ : std_logic;
SIGNAL \RegFile[2][17]~q\ : std_logic;
SIGNAL \RegFile[4][17]~feeder_combout\ : std_logic;
SIGNAL \RegFile[4][17]~q\ : std_logic;
SIGNAL \RegFile[6][17]~feeder_combout\ : std_logic;
SIGNAL \RegFile[6][17]~q\ : std_logic;
SIGNAL \RegFile[5][17]~q\ : std_logic;
SIGNAL \RegFile[7][17]~q\ : std_logic;
SIGNAL \Mux73~0_combout\ : std_logic;
SIGNAL \RegFile[1][17]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux73~26_combout\ : std_logic;
SIGNAL \RegFile[31][17]~q\ : std_logic;
SIGNAL \RegFile[30][17]~q\ : std_logic;
SIGNAL \RegFile[29][17]~q\ : std_logic;
SIGNAL \RegFile[25][17]~q\ : std_logic;
SIGNAL \RegFile[27][17]~q\ : std_logic;
SIGNAL \RegFile[26][17]~feeder_combout\ : std_logic;
SIGNAL \RegFile[26][17]~q\ : std_logic;
SIGNAL \RegFile[24][17]~q\ : std_logic;
SIGNAL \Mux73~22_combout\ : std_logic;
SIGNAL \RegFile[28][17]~feeder_combout\ : std_logic;
SIGNAL \RegFile[28][17]~q\ : std_logic;
SIGNAL \Mux73~9_combout\ : std_logic;
SIGNAL \RegFile[21][17]~feeder_combout\ : std_logic;
SIGNAL \RegFile[21][17]~q\ : std_logic;
SIGNAL \RegFile[23][17]~q\ : std_logic;
SIGNAL \RegFile[22][17]~feeder_combout\ : std_logic;
SIGNAL \RegFile[22][17]~q\ : std_logic;
SIGNAL \RegFile[17][17]~q\ : std_logic;
SIGNAL \RegFile[19][17]~q\ : std_logic;
SIGNAL \RegFile[18][17]~feeder_combout\ : std_logic;
SIGNAL \RegFile[18][17]~q\ : std_logic;
SIGNAL \RegFile[16][17]~feeder_combout\ : std_logic;
SIGNAL \RegFile[16][17]~q\ : std_logic;
SIGNAL \Mux73~18_combout\ : std_logic;
SIGNAL \RegFile[20][17]~q\ : std_logic;
SIGNAL \Mux73~5_combout\ : std_logic;
SIGNAL \RegFile[15][17]~q\ : std_logic;
SIGNAL \RegFile[14][17]~feeder_combout\ : std_logic;
SIGNAL \RegFile[14][17]~q\ : std_logic;
SIGNAL \RegFile[11][17]~q\ : std_logic;
SIGNAL \RegFile[9][17]~q\ : std_logic;
SIGNAL \RegFile[10][17]~feeder_combout\ : std_logic;
SIGNAL \RegFile[10][17]~q\ : std_logic;
SIGNAL \RegFile[8][17]~q\ : std_logic;
SIGNAL \Mux73~14_combout\ : std_logic;
SIGNAL \RegFile[12][17]~q\ : std_logic;
SIGNAL \Mux73~1_combout\ : std_logic;
SIGNAL \Mux73~13_combout\ : std_logic;
SIGNAL \Mux237~0_combout\ : std_logic;
SIGNAL \ShiftRight1~10_combout\ : std_logic;
SIGNAL \ShiftRight1~10_OTERM265\ : std_logic;
SIGNAL \ShiftRight1~42_combout\ : std_logic;
SIGNAL \Selector27~4_combout\ : std_logic;
SIGNAL \Add2~17_OTERM727_OTERM841\ : std_logic;
SIGNAL \Add1~6\ : std_logic;
SIGNAL \Add1~10\ : std_logic;
SIGNAL \Add1~14\ : std_logic;
SIGNAL \Add1~18\ : std_logic;
SIGNAL \Add1~21_sumout\ : std_logic;
SIGNAL \Add2~6\ : std_logic;
SIGNAL \Add2~7\ : std_logic;
SIGNAL \Add2~10\ : std_logic;
SIGNAL \Add2~11\ : std_logic;
SIGNAL \Add2~14\ : std_logic;
SIGNAL \Add2~15\ : std_logic;
SIGNAL \Add2~18\ : std_logic;
SIGNAL \Add2~19\ : std_logic;
SIGNAL \Add2~21_sumout\ : std_logic;
SIGNAL \Selector27~1_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[5]~0_RESYN1092_BDD1093\ : std_logic;
SIGNAL \Comb:vRegWriteData[5]~0_combout\ : std_logic;
SIGNAL \Selector16~0_combout\ : std_logic;
SIGNAL \Selector16~0_OTERM393\ : std_logic;
SIGNAL \Mux135~0_combout\ : std_logic;
SIGNAL \RegFile[23][19]~q\ : std_logic;
SIGNAL \RegFile[21][19]~q\ : std_logic;
SIGNAL \RegFile[22][19]~feeder_combout\ : std_logic;
SIGNAL \RegFile[22][19]~q\ : std_logic;
SIGNAL \RegFile[19][19]~q\ : std_logic;
SIGNAL \RegFile[17][19]~q\ : std_logic;
SIGNAL \RegFile[18][19]~feeder_combout\ : std_logic;
SIGNAL \RegFile[18][19]~q\ : std_logic;
SIGNAL \RegFile[16][19]~q\ : std_logic;
SIGNAL \Mux103~18_combout\ : std_logic;
SIGNAL \RegFile[20][19]~q\ : std_logic;
SIGNAL \Mux103~5_combout\ : std_logic;
SIGNAL \RegFile[2][19]~q\ : std_logic;
SIGNAL \RegFile[7][19]~q\ : std_logic;
SIGNAL \RegFile[6][19]~feeder_combout\ : std_logic;
SIGNAL \RegFile[6][19]~q\ : std_logic;
SIGNAL \RegFile[4][19]~q\ : std_logic;
SIGNAL \RegFile[5][19]~q\ : std_logic;
SIGNAL \Mux103~0_combout\ : std_logic;
SIGNAL \RegFile[1][19]~feeder_combout\ : std_logic;
SIGNAL \RegFile[1][19]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux103~26_combout\ : std_logic;
SIGNAL \RegFile[29][19]~q\ : std_logic;
SIGNAL \RegFile[30][19]~q\ : std_logic;
SIGNAL \RegFile[31][19]~q\ : std_logic;
SIGNAL \RegFile[25][19]~q\ : std_logic;
SIGNAL \RegFile[27][19]~q\ : std_logic;
SIGNAL \RegFile[26][19]~feeder_combout\ : std_logic;
SIGNAL \RegFile[26][19]~q\ : std_logic;
SIGNAL \RegFile[24][19]~q\ : std_logic;
SIGNAL \Mux103~22_combout\ : std_logic;
SIGNAL \RegFile[28][19]~q\ : std_logic;
SIGNAL \Mux103~9_combout\ : std_logic;
SIGNAL \RegFile[13][19]~q\ : std_logic;
SIGNAL \RegFile[15][19]~q\ : std_logic;
SIGNAL \RegFile[14][19]~q\ : std_logic;
SIGNAL \RegFile[9][19]~q\ : std_logic;
SIGNAL \RegFile[10][19]~feeder_combout\ : std_logic;
SIGNAL \RegFile[10][19]~q\ : std_logic;
SIGNAL \RegFile[11][19]~feeder_combout\ : std_logic;
SIGNAL \RegFile[11][19]~q\ : std_logic;
SIGNAL \RegFile[8][19]~q\ : std_logic;
SIGNAL \Mux103~14_combout\ : std_logic;
SIGNAL \RegFile[12][19]~q\ : std_logic;
SIGNAL \Mux103~1_combout\ : std_logic;
SIGNAL \Mux103~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[19]~2_combout\ : std_logic;
SIGNAL \Selector13~4_combout\ : std_logic;
SIGNAL \Selector13~5_combout\ : std_logic;
SIGNAL \Mux136~0_combout\ : std_logic;
SIGNAL \RegFile[15][18]~q\ : std_logic;
SIGNAL \RegFile[13][18]~q\ : std_logic;
SIGNAL \RegFile[14][18]~feeder_combout\ : std_logic;
SIGNAL \RegFile[14][18]~q\ : std_logic;
SIGNAL \RegFile[9][18]~q\ : std_logic;
SIGNAL \RegFile[10][18]~feeder_combout\ : std_logic;
SIGNAL \RegFile[10][18]~DUPLICATE_q\ : std_logic;
SIGNAL \RegFile[11][18]~q\ : std_logic;
SIGNAL \RegFile[8][18]~feeder_combout\ : std_logic;
SIGNAL \RegFile[8][18]~q\ : std_logic;
SIGNAL \Mux104~14_combout\ : std_logic;
SIGNAL \RegFile[12][18]~q\ : std_logic;
SIGNAL \Mux104~1_combout\ : std_logic;
SIGNAL \RegFile[23][18]~q\ : std_logic;
SIGNAL \RegFile[22][18]~feeder_combout\ : std_logic;
SIGNAL \RegFile[22][18]~q\ : std_logic;
SIGNAL \RegFile[19][18]~q\ : std_logic;
SIGNAL \RegFile[18][18]~q\ : std_logic;
SIGNAL \RegFile[17][18]~q\ : std_logic;
SIGNAL \RegFile[16][18]~q\ : std_logic;
SIGNAL \Mux104~18_combout\ : std_logic;
SIGNAL \RegFile[20][18]~feeder_combout\ : std_logic;
SIGNAL \RegFile[20][18]~q\ : std_logic;
SIGNAL \Mux104~5_combout\ : std_logic;
SIGNAL \RegFile[3][18]~q\ : std_logic;
SIGNAL \RegFile[2][18]~q\ : std_logic;
SIGNAL \RegFile[5][18]~q\ : std_logic;
SIGNAL \RegFile[4][18]~DUPLICATE_q\ : std_logic;
SIGNAL \RegFile[6][18]~feeder_combout\ : std_logic;
SIGNAL \RegFile[6][18]~DUPLICATE_q\ : std_logic;
SIGNAL \RegFile[7][18]~q\ : std_logic;
SIGNAL \Mux104~0_combout\ : std_logic;
SIGNAL \RegFile[1][18]~feeder_combout\ : std_logic;
SIGNAL \RegFile[1][18]~q\ : std_logic;
SIGNAL \Mux104~26_combout\ : std_logic;
SIGNAL \RegFile[29][18]~q\ : std_logic;
SIGNAL \RegFile[30][18]~feeder_combout\ : std_logic;
SIGNAL \RegFile[30][18]~q\ : std_logic;
SIGNAL \RegFile[31][18]~q\ : std_logic;
SIGNAL \RegFile[25][18]~q\ : std_logic;
SIGNAL \RegFile[26][18]~feeder_combout\ : std_logic;
SIGNAL \RegFile[26][18]~q\ : std_logic;
SIGNAL \RegFile[27][18]~q\ : std_logic;
SIGNAL \RegFile[24][18]~feeder_combout\ : std_logic;
SIGNAL \RegFile[24][18]~q\ : std_logic;
SIGNAL \Mux104~22_combout\ : std_logic;
SIGNAL \RegFile[28][18]~feeder_combout\ : std_logic;
SIGNAL \RegFile[28][18]~q\ : std_logic;
SIGNAL \Mux104~9_combout\ : std_logic;
SIGNAL \Mux104~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[18]~3_combout\ : std_logic;
SIGNAL \Add2~65_OTERM703_OTERM805\ : std_logic;
SIGNAL \Mux138~0_combout\ : std_logic;
SIGNAL \Add0~57_sumout\ : std_logic;
SIGNAL \R.regWriteData[16]~feeder_combout\ : std_logic;
SIGNAL \Add2~65_OTERM703_OTERM809\ : std_logic;
SIGNAL \Add1~58\ : std_logic;
SIGNAL \Add1~62\ : std_logic;
SIGNAL \Add1~65_sumout\ : std_logic;
SIGNAL \Add2~25_OTERM723_OTERM833\ : std_logic;
SIGNAL \Add2~22\ : std_logic;
SIGNAL \Add2~23\ : std_logic;
SIGNAL \Add2~26\ : std_logic;
SIGNAL \Add2~27\ : std_logic;
SIGNAL \Add2~30\ : std_logic;
SIGNAL \Add2~31\ : std_logic;
SIGNAL \Add2~34\ : std_logic;
SIGNAL \Add2~35\ : std_logic;
SIGNAL \Add2~38\ : std_logic;
SIGNAL \Add2~39\ : std_logic;
SIGNAL \Add2~42\ : std_logic;
SIGNAL \Add2~43\ : std_logic;
SIGNAL \Add2~46\ : std_logic;
SIGNAL \Add2~47\ : std_logic;
SIGNAL \Add2~50\ : std_logic;
SIGNAL \Add2~51\ : std_logic;
SIGNAL \Add2~54\ : std_logic;
SIGNAL \Add2~55\ : std_logic;
SIGNAL \Add2~59\ : std_logic;
SIGNAL \Add2~62\ : std_logic;
SIGNAL \Add2~63\ : std_logic;
SIGNAL \Add2~65_sumout\ : std_logic;
SIGNAL \Comb:vRegWriteData[24]~1_combout\ : std_logic;
SIGNAL \avm_d_readdata[23]~input_o\ : std_logic;
SIGNAL \avm_d_readdata[31]~input_o\ : std_logic;
SIGNAL \avm_d_readdata[8]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[16]~0_RESYN1724_BDD1725\ : std_logic;
SIGNAL \Comb:vRegWriteData[16]~0_RESYN1726_BDD1727\ : std_logic;
SIGNAL \Comb:vRegWriteData[16]~0_RESYN1728_BDD1729\ : std_logic;
SIGNAL \Comb:vRegWriteData[16]~0_combout\ : std_logic;
SIGNAL \RegFile[23][16]~q\ : std_logic;
SIGNAL \RegFile[21][16]~q\ : std_logic;
SIGNAL \RegFile[22][16]~q\ : std_logic;
SIGNAL \RegFile[19][16]~q\ : std_logic;
SIGNAL \RegFile[18][16]~q\ : std_logic;
SIGNAL \RegFile[17][16]~q\ : std_logic;
SIGNAL \RegFile[16][16]~q\ : std_logic;
SIGNAL \Mux106~18_combout\ : std_logic;
SIGNAL \RegFile[20][16]~q\ : std_logic;
SIGNAL \Mux106~5_combout\ : std_logic;
SIGNAL \RegFile[15][16]~q\ : std_logic;
SIGNAL \RegFile[14][16]~DUPLICATE_q\ : std_logic;
SIGNAL \RegFile[13][16]~q\ : std_logic;
SIGNAL \RegFile[9][16]~q\ : std_logic;
SIGNAL \RegFile[10][16]~feeder_combout\ : std_logic;
SIGNAL \RegFile[10][16]~q\ : std_logic;
SIGNAL \RegFile[11][16]~q\ : std_logic;
SIGNAL \RegFile[8][16]~feeder_combout\ : std_logic;
SIGNAL \RegFile[8][16]~q\ : std_logic;
SIGNAL \Mux106~14_combout\ : std_logic;
SIGNAL \RegFile[12][16]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux106~1_combout\ : std_logic;
SIGNAL \RegFile[3][16]~q\ : std_logic;
SIGNAL \RegFile[2][16]~q\ : std_logic;
SIGNAL \RegFile[4][16]~feeder_combout\ : std_logic;
SIGNAL \RegFile[4][16]~q\ : std_logic;
SIGNAL \RegFile[5][16]~DUPLICATE_q\ : std_logic;
SIGNAL \RegFile[7][16]~q\ : std_logic;
SIGNAL \RegFile[6][16]~q\ : std_logic;
SIGNAL \Mux106~0_combout\ : std_logic;
SIGNAL \RegFile[1][16]~q\ : std_logic;
SIGNAL \Mux106~26_combout\ : std_logic;
SIGNAL \RegFile[31][16]~q\ : std_logic;
SIGNAL \RegFile[30][16]~feeder_combout\ : std_logic;
SIGNAL \RegFile[30][16]~q\ : std_logic;
SIGNAL \RegFile[29][16]~q\ : std_logic;
SIGNAL \RegFile[25][16]~q\ : std_logic;
SIGNAL \RegFile[26][16]~feeder_combout\ : std_logic;
SIGNAL \RegFile[26][16]~q\ : std_logic;
SIGNAL \RegFile[27][16]~q\ : std_logic;
SIGNAL \RegFile[24][16]~feeder_combout\ : std_logic;
SIGNAL \RegFile[24][16]~q\ : std_logic;
SIGNAL \Mux106~22_combout\ : std_logic;
SIGNAL \RegFile[28][16]~feeder_combout\ : std_logic;
SIGNAL \RegFile[28][16]~q\ : std_logic;
SIGNAL \Mux106~9_combout\ : std_logic;
SIGNAL \Mux106~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[16]~5_combout\ : std_logic;
SIGNAL \Add2~65_OTERM703_OTERM811\ : std_logic;
SIGNAL \Add1~66\ : std_logic;
SIGNAL \Add1~70\ : std_logic;
SIGNAL \Add1~74\ : std_logic;
SIGNAL \Add1~77_sumout\ : std_logic;
SIGNAL \Add2~66\ : std_logic;
SIGNAL \Add2~67\ : std_logic;
SIGNAL \Add2~70\ : std_logic;
SIGNAL \Add2~71\ : std_logic;
SIGNAL \Add2~74\ : std_logic;
SIGNAL \Add2~75\ : std_logic;
SIGNAL \Add2~77_sumout\ : std_logic;
SIGNAL \Selector13~1_combout\ : std_logic;
SIGNAL \Add2~79\ : std_logic;
SIGNAL \Add2~83\ : std_logic;
SIGNAL \Add2~85_sumout\ : std_logic;
SIGNAL \Selector13~3_combout\ : std_logic;
SIGNAL \Selector11~0_combout\ : std_logic;
SIGNAL \ShiftLeft0~12_combout\ : std_logic;
SIGNAL \ShiftLeft0~12_OTERM791\ : std_logic;
SIGNAL \ShiftLeft0~26_combout\ : std_logic;
SIGNAL \ShiftLeft0~26_OTERM739\ : std_logic;
SIGNAL \ShiftLeft0~18_combout\ : std_logic;
SIGNAL \ShiftLeft0~18_OTERM289\ : std_logic;
SIGNAL \ShiftLeft0~34_combout\ : std_logic;
SIGNAL \ShiftLeft0~34_OTERM299\ : std_logic;
SIGNAL \ShiftLeft0~35_combout\ : std_logic;
SIGNAL \Selector11~1_combout\ : std_logic;
SIGNAL \Add1~78\ : std_logic;
SIGNAL \Add1~82\ : std_logic;
SIGNAL \Add1~85_sumout\ : std_logic;
SIGNAL \Equal3~5_RESYN1100_BDD1101\ : std_logic;
SIGNAL \Equal3~5_RESYN1102_BDD1103\ : std_logic;
SIGNAL \Equal3~5_combout\ : std_logic;
SIGNAL \R.statusReg[0]_OTERM9_OTERM473\ : std_logic;
SIGNAL \Add2~87\ : std_logic;
SIGNAL \Add2~91\ : std_logic;
SIGNAL \Add2~95\ : std_logic;
SIGNAL \Add2~99\ : std_logic;
SIGNAL \Add2~103\ : std_logic;
SIGNAL \Add2~107\ : std_logic;
SIGNAL \Add2~109_sumout\ : std_logic;
SIGNAL \ShiftLeft0~38_combout\ : std_logic;
SIGNAL \ShiftLeft0~38_OTERM789\ : std_logic;
SIGNAL \ShiftLeft0~47_combout\ : std_logic;
SIGNAL \ShiftLeft0~47_OTERM759\ : std_logic;
SIGNAL \ShiftLeft0~30_combout\ : std_logic;
SIGNAL \ShiftLeft0~30_OTERM601\ : std_logic;
SIGNAL \ShiftLeft0~22_combout\ : std_logic;
SIGNAL \ShiftLeft0~22_OTERM737\ : std_logic;
SIGNAL \ShiftLeft0~48_combout\ : std_logic;
SIGNAL \ShiftRight1~32_combout\ : std_logic;
SIGNAL \ShiftRight1~32_OTERM21\ : std_logic;
SIGNAL \ShiftRight0~4_combout\ : std_logic;
SIGNAL \ShiftRight0~4_OTERM31\ : std_logic;
SIGNAL \Selector5~0_combout\ : std_logic;
SIGNAL \Selector5~1_combout\ : std_logic;
SIGNAL \Selector5~2_combout\ : std_logic;
SIGNAL \ShiftLeft0~9_combout\ : std_logic;
SIGNAL \ShiftLeft0~9_OTERM461\ : std_logic;
SIGNAL \ShiftLeft0~15_combout\ : std_logic;
SIGNAL \Selector5~3_combout\ : std_logic;
SIGNAL \Selector5~4_combout\ : std_logic;
SIGNAL \Selector5~5_combout\ : std_logic;
SIGNAL \vAluRes~35_combout\ : std_logic;
SIGNAL \vAluRes~24_combout\ : std_logic;
SIGNAL \R.statusReg[0]_OTERM9_OTERM467\ : std_logic;
SIGNAL \Add1~69_sumout\ : std_logic;
SIGNAL \Equal3~14_combout\ : std_logic;
SIGNAL \ShiftLeft0~1_combout\ : std_logic;
SIGNAL \ShiftLeft0~1_OTERM255\ : std_logic;
SIGNAL \Selector15~2_RTM0743_combout\ : std_logic;
SIGNAL \Selector15~2_OTERM741\ : std_logic;
SIGNAL \Selector15~3_combout\ : std_logic;
SIGNAL \ShiftLeft0~27_combout\ : std_logic;
SIGNAL \Selector15~4_combout\ : std_logic;
SIGNAL \ShiftRight1~14_combout\ : std_logic;
SIGNAL \Selector15~0_combout\ : std_logic;
SIGNAL \Equal3~15_combout\ : std_logic;
SIGNAL \Equal3~4_combout\ : std_logic;
SIGNAL \R.statusReg[0]_OTERM9_OTERM471\ : std_logic;
SIGNAL \R.statusReg[0]_OTERM9_OTERM463\ : std_logic;
SIGNAL \ShiftLeft0~0_combout\ : std_logic;
SIGNAL \ShiftLeft0~0_OTERM263\ : std_logic;
SIGNAL \ShiftLeft0~16_combout\ : std_logic;
SIGNAL \ShiftLeft0~16_OTERM287\ : std_logic;
SIGNAL \ShiftLeft0~17_combout\ : std_logic;
SIGNAL \Selector20~2_combout\ : std_logic;
SIGNAL \Selector20~0_combout\ : std_logic;
SIGNAL \Selector20~0_OTERM769\ : std_logic;
SIGNAL \ShiftRight1~3_combout\ : std_logic;
SIGNAL \ShiftRight1~3_OTERM13\ : std_logic;
SIGNAL \Selector20~1_combout\ : std_logic;
SIGNAL \ShiftRight1~0_combout\ : std_logic;
SIGNAL \ShiftRight1~0_OTERM257\ : std_logic;
SIGNAL \ShiftRight1~8_combout\ : std_logic;
SIGNAL \ShiftRight1~8_OTERM261\ : std_logic;
SIGNAL \ShiftRight1~1_combout\ : std_logic;
SIGNAL \ShiftRight1~1_OTERM33\ : std_logic;
SIGNAL \ShiftRight1~2_combout\ : std_logic;
SIGNAL \ShiftRight1~2_OTERM49\ : std_logic;
SIGNAL \ShiftRight1~51_combout\ : std_logic;
SIGNAL \Selector20~3_combout\ : std_logic;
SIGNAL \ShiftRight1~31_combout\ : std_logic;
SIGNAL \ShiftRight1~31_OTERM45\ : std_logic;
SIGNAL \Selector25~2_combout\ : std_logic;
SIGNAL \ShiftRight1~30_combout\ : std_logic;
SIGNAL \ShiftRight1~30_OTERM39\ : std_logic;
SIGNAL \ShiftRight1~37_combout\ : std_logic;
SIGNAL \ShiftRight1~37_OTERM283\ : std_logic;
SIGNAL \ShiftRight1~35_combout\ : std_logic;
SIGNAL \ShiftRight1~35_OTERM279\ : std_logic;
SIGNAL \ShiftRight1~45_combout\ : std_logic;
SIGNAL \Selector25~3_RTM0799_combout\ : std_logic;
SIGNAL \Selector25~3_OTERM797\ : std_logic;
SIGNAL \Selector25~4_combout\ : std_logic;
SIGNAL \Selector25~6_RESYN1116_BDD1117\ : std_logic;
SIGNAL \Selector25~1_combout\ : std_logic;
SIGNAL \Add2~29_sumout\ : std_logic;
SIGNAL \Selector25~6_combout\ : std_logic;
SIGNAL \Add1~49_sumout\ : std_logic;
SIGNAL \Selector20~6_combout\ : std_logic;
SIGNAL \Equal3~10_combout\ : std_logic;
SIGNAL \Equal3~3_combout\ : std_logic;
SIGNAL \R.statusReg[0]_OTERM9_OTERM469\ : std_logic;
SIGNAL \LessThan1~31_combout\ : std_logic;
SIGNAL \Selector10~2_combout\ : std_logic;
SIGNAL \Selector10~3_combout\ : std_logic;
SIGNAL \Selector10~4_combout\ : std_logic;
SIGNAL \ShiftLeft0~20_combout\ : std_logic;
SIGNAL \ShiftLeft0~20_OTERM291\ : std_logic;
SIGNAL \ShiftLeft0~13_combout\ : std_logic;
SIGNAL \ShiftLeft0~13_OTERM285\ : std_logic;
SIGNAL \ShiftLeft0~28_combout\ : std_logic;
SIGNAL \ShiftLeft0~28_OTERM295\ : std_logic;
SIGNAL \ShiftLeft0~37_combout\ : std_logic;
SIGNAL \ShiftRight0~2_combout\ : std_logic;
SIGNAL \ShiftRight0~2_OTERM25\ : std_logic;
SIGNAL \Selector10~0_combout\ : std_logic;
SIGNAL \Selector10~1_combout\ : std_logic;
SIGNAL \Add2~89_sumout\ : std_logic;
SIGNAL \Selector10~5_combout\ : std_logic;
SIGNAL \vAluRes~34_combout\ : std_logic;
SIGNAL \vAluRes~19_combout\ : std_logic;
SIGNAL \R.statusReg[0]_OTERM9_OTERM465\ : std_logic;
SIGNAL \Equal3~6_combout\ : std_logic;
SIGNAL \ShiftLeft0~32_combout\ : std_logic;
SIGNAL \ShiftLeft0~32_OTERM297\ : std_logic;
SIGNAL \ShiftLeft0~40_combout\ : std_logic;
SIGNAL \ShiftLeft0~40_OTERM755\ : std_logic;
SIGNAL \ShiftLeft0~49_combout\ : std_logic;
SIGNAL \ShiftLeft0~49_OTERM761\ : std_logic;
SIGNAL \ShiftLeft0~50_combout\ : std_logic;
SIGNAL \Selector4~0_combout\ : std_logic;
SIGNAL \Selector20~5_combout\ : std_logic;
SIGNAL \Selector4~1_combout\ : std_logic;
SIGNAL \Add2~111\ : std_logic;
SIGNAL \Add2~113_sumout\ : std_logic;
SIGNAL \Selector4~2_combout\ : std_logic;
SIGNAL \vAluRes~48_combout\ : std_logic;
SIGNAL \R.statusReg[0]_OTERM5\ : std_logic;
SIGNAL \R.statusReg[0]_OTERM7_OTERM491\ : std_logic;
SIGNAL \ShiftLeft0~23_combout\ : std_logic;
SIGNAL \Selector1~0_RTM0773_combout\ : std_logic;
SIGNAL \Selector1~0_OTERM771\ : std_logic;
SIGNAL \Selector1~1_combout\ : std_logic;
SIGNAL \ShiftLeft0~55_combout\ : std_logic;
SIGNAL \ShiftLeft0~55_OTERM767\ : std_logic;
SIGNAL \ShiftLeft0~56_combout\ : std_logic;
SIGNAL \Selector1~2_combout\ : std_logic;
SIGNAL \R.statusReg[0]_OTERM7_OTERM481\ : std_logic;
SIGNAL \R.statusReg[0]_OTERM7_OTERM483\ : std_logic;
SIGNAL \Equal3~19_combout\ : std_logic;
SIGNAL \R.statusReg[0]_OTERM7_OTERM489\ : std_logic;
SIGNAL \Add1~122\ : std_logic;
SIGNAL \Add1~125_sumout\ : std_logic;
SIGNAL \Add2~101_sumout\ : std_logic;
SIGNAL \Add1~94\ : std_logic;
SIGNAL \Add1~98\ : std_logic;
SIGNAL \Add1~101_sumout\ : std_logic;
SIGNAL \Selector7~3_combout\ : std_logic;
SIGNAL \vAluRes~26_combout\ : std_logic;
SIGNAL \Equal3~18_combout\ : std_logic;
SIGNAL \R.statusReg[0]_OTERM7_OTERM487\ : std_logic;
SIGNAL \Add1~105_sumout\ : std_logic;
SIGNAL \Add2~105_sumout\ : std_logic;
SIGNAL \vAluRes~27_combout\ : std_logic;
SIGNAL \R.statusReg[0]_OTERM7_OTERM485\ : std_logic;
SIGNAL \Equal3~2_combout\ : std_logic;
SIGNAL \vAluRes~33_combout\ : std_logic;
SIGNAL \Add1~81_sumout\ : std_logic;
SIGNAL \vAluRes~17_combout\ : std_logic;
SIGNAL \R.aluRes[0]~DUPLICATE_q\ : std_logic;
SIGNAL \vAluRes~0_combout\ : std_logic;
SIGNAL \Equal3~1_combout\ : std_logic;
SIGNAL \R.statusReg[0]_OTERM11_OTERM375\ : std_logic;
SIGNAL \R.statusReg[0]_OTERM11_OTERM371\ : std_logic;
SIGNAL \R.statusReg[0]_OTERM11_OTERM369\ : std_logic;
SIGNAL \R.statusReg[0]_OTERM11_OTERM373\ : std_logic;
SIGNAL \R.statusReg[0]_OTERM11_OTERM367\ : std_logic;
SIGNAL \Add2~57_sumout\ : std_logic;
SIGNAL \Selector23~1_combout\ : std_logic;
SIGNAL \Add2~37_sumout\ : std_logic;
SIGNAL \Selector23~2_combout\ : std_logic;
SIGNAL \Selector23~3_RTM0425_combout\ : std_logic;
SIGNAL \Selector23~3_OTERM423\ : std_logic;
SIGNAL \Selector23~4_combout\ : std_logic;
SIGNAL \Selector23~7_combout\ : std_logic;
SIGNAL \Selector23~6_combout\ : std_logic;
SIGNAL \Selector18~5_combout\ : std_logic;
SIGNAL \Equal3~11_combout\ : std_logic;
SIGNAL \Equal3~7_combout\ : std_logic;
SIGNAL \R.statusReg[0]_OTERM11_OTERM377_OTERM595\ : std_logic;
SIGNAL \R.statusReg[0]_OTERM11_OTERM377_OTERM593\ : std_logic;
SIGNAL \ShiftLeft0~29_combout\ : std_logic;
SIGNAL \ShiftRight1~25_combout\ : std_logic;
SIGNAL \ShiftRight1~25_OTERM277\ : std_logic;
SIGNAL \ShiftRight0~3_combout\ : std_logic;
SIGNAL \Selector14~0_combout\ : std_logic;
SIGNAL \Selector14~5_combout\ : std_logic;
SIGNAL \Selector14~4_combout\ : std_logic;
SIGNAL \Equal3~12_RESYN1054_BDD1055\ : std_logic;
SIGNAL \Equal3~12_combout\ : std_logic;
SIGNAL \R.statusReg[0]_OTERM11_OTERM377_OTERM597\ : std_logic;
SIGNAL \Equal3~13_combout\ : std_logic;
SIGNAL \Equal3~9_combout\ : std_logic;
SIGNAL \R.aluRes[30]~DUPLICATE_q\ : std_logic;
SIGNAL \vAluRes~40_combout\ : std_logic;
SIGNAL \R.statusReg[0]_OTERM1\ : std_logic;
SIGNAL \Add2~115\ : std_logic;
SIGNAL \Add2~117_sumout\ : std_logic;
SIGNAL \vAluRes~44_combout\ : std_logic;
SIGNAL \R.statusReg[0]_OTERM3\ : std_logic;
SIGNAL \Equal3~8_combout\ : std_logic;
SIGNAL \vAluRes~36_combout\ : std_logic;
SIGNAL \ShiftLeft0~57_combout\ : std_logic;
SIGNAL \ShiftLeft0~58_combout\ : std_logic;
SIGNAL \Selector0~0_combout\ : std_logic;
SIGNAL \Add1~126\ : std_logic;
SIGNAL \Add1~129_sumout\ : std_logic;
SIGNAL \Add2~119\ : std_logic;
SIGNAL \Add2~122\ : std_logic;
SIGNAL \Add2~123\ : std_logic;
SIGNAL \Add2~126\ : std_logic;
SIGNAL \Add2~127\ : std_logic;
SIGNAL \Add2~129_sumout\ : std_logic;
SIGNAL \Selector0~1_combout\ : std_logic;
SIGNAL \Mux58~0_combout\ : std_logic;
SIGNAL \NxR~8_combout\ : std_logic;
SIGNAL \R.jumpToAdr~q\ : std_logic;
SIGNAL \RegFile[29][5]~q\ : std_logic;
SIGNAL \Mux85~22_combout\ : std_logic;
SIGNAL \Mux85~9_combout\ : std_logic;
SIGNAL \Mux85~14_combout\ : std_logic;
SIGNAL \Mux85~1_combout\ : std_logic;
SIGNAL \Mux85~0_combout\ : std_logic;
SIGNAL \Mux85~26_combout\ : std_logic;
SIGNAL \RegFile[16][5]~q\ : std_logic;
SIGNAL \Mux85~18_combout\ : std_logic;
SIGNAL \Mux85~5_combout\ : std_logic;
SIGNAL \Mux85~13_combout\ : std_logic;
SIGNAL \Mux249~0_combout\ : std_logic;
SIGNAL \ShiftLeft0~8_combout\ : std_logic;
SIGNAL \ShiftLeft0~8_OTERM207\ : std_logic;
SIGNAL \Selector26~1_combout\ : std_logic;
SIGNAL \ShiftRight0~9_combout\ : std_logic;
SIGNAL \ShiftRight1~22_combout\ : std_logic;
SIGNAL \ShiftRight1~22_OTERM273\ : std_logic;
SIGNAL \ShiftRight1~23_combout\ : std_logic;
SIGNAL \ShiftRight1~23_OTERM275\ : std_logic;
SIGNAL \ShiftRight1~21_combout\ : std_logic;
SIGNAL \ShiftRight1~21_OTERM271\ : std_logic;
SIGNAL \ShiftRight1~44_combout\ : std_logic;
SIGNAL \Selector26~3_combout\ : std_logic;
SIGNAL \Add2~25_sumout\ : std_logic;
SIGNAL \Add1~22\ : std_logic;
SIGNAL \Add1~25_sumout\ : std_logic;
SIGNAL \Selector26~0_combout\ : std_logic;
SIGNAL \avm_d_readdata[30]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[6]~0_RESYN1098_BDD1099\ : std_logic;
SIGNAL \Comb:vRegWriteData[6]~0_combout\ : std_logic;
SIGNAL \RegFile[21][6]~q\ : std_logic;
SIGNAL \RegFile[23][6]~q\ : std_logic;
SIGNAL \RegFile[22][6]~q\ : std_logic;
SIGNAL \RegFile[17][6]~q\ : std_logic;
SIGNAL \RegFile[18][6]~feeder_combout\ : std_logic;
SIGNAL \RegFile[18][6]~q\ : std_logic;
SIGNAL \RegFile[19][6]~q\ : std_logic;
SIGNAL \RegFile[16][6]~feeder_combout\ : std_logic;
SIGNAL \RegFile[16][6]~q\ : std_logic;
SIGNAL \Mux116~18_combout\ : std_logic;
SIGNAL \RegFile[20][6]~q\ : std_logic;
SIGNAL \Mux116~5_combout\ : std_logic;
SIGNAL \RegFile[3][6]~q\ : std_logic;
SIGNAL \RegFile[2][6]~q\ : std_logic;
SIGNAL \RegFile[4][6]~q\ : std_logic;
SIGNAL \RegFile[5][6]~q\ : std_logic;
SIGNAL \RegFile[7][6]~q\ : std_logic;
SIGNAL \RegFile[6][6]~q\ : std_logic;
SIGNAL \Mux116~0_combout\ : std_logic;
SIGNAL \RegFile[1][6]~q\ : std_logic;
SIGNAL \Mux116~26_combout\ : std_logic;
SIGNAL \RegFile[31][6]~feeder_combout\ : std_logic;
SIGNAL \RegFile[31][6]~q\ : std_logic;
SIGNAL \RegFile[30][6]~feeder_combout\ : std_logic;
SIGNAL \RegFile[30][6]~q\ : std_logic;
SIGNAL \RegFile[29][6]~q\ : std_logic;
SIGNAL \RegFile[27][6]~feeder_combout\ : std_logic;
SIGNAL \RegFile[27][6]~q\ : std_logic;
SIGNAL \RegFile[25][6]~q\ : std_logic;
SIGNAL \RegFile[26][6]~feeder_combout\ : std_logic;
SIGNAL \RegFile[26][6]~q\ : std_logic;
SIGNAL \RegFile[24][6]~feeder_combout\ : std_logic;
SIGNAL \RegFile[24][6]~q\ : std_logic;
SIGNAL \Mux116~22_combout\ : std_logic;
SIGNAL \RegFile[28][6]~q\ : std_logic;
SIGNAL \Mux116~9_combout\ : std_logic;
SIGNAL \RegFile[13][6]~q\ : std_logic;
SIGNAL \RegFile[15][6]~q\ : std_logic;
SIGNAL \RegFile[14][6]~q\ : std_logic;
SIGNAL \RegFile[9][6]~q\ : std_logic;
SIGNAL \RegFile[10][6]~feeder_combout\ : std_logic;
SIGNAL \RegFile[10][6]~q\ : std_logic;
SIGNAL \RegFile[11][6]~q\ : std_logic;
SIGNAL \RegFile[8][6]~q\ : std_logic;
SIGNAL \Mux116~14_combout\ : std_logic;
SIGNAL \RegFile[12][6]~feeder_combout\ : std_logic;
SIGNAL \RegFile[12][6]~q\ : std_logic;
SIGNAL \Mux116~1_combout\ : std_logic;
SIGNAL \Mux116~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[6]~15_combout\ : std_logic;
SIGNAL \Add2~25_OTERM723_OTERM835\ : std_logic;
SIGNAL \Add1~26\ : std_logic;
SIGNAL \Add1~30\ : std_logic;
SIGNAL \Add1~34\ : std_logic;
SIGNAL \Add1~37_sumout\ : std_logic;
SIGNAL \Comb:vRegWriteData[9]~1_RESYN1080_BDD1081\ : std_logic;
SIGNAL \avm_d_readdata[17]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[9]~1_RESYN1078_BDD1079\ : std_logic;
SIGNAL \Comb:vRegWriteData[9]~1_combout\ : std_logic;
SIGNAL \RegFile[13][9]~q\ : std_logic;
SIGNAL \RegFile[14][9]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux113~14_combout\ : std_logic;
SIGNAL \Mux113~1_combout\ : std_logic;
SIGNAL \Mux113~22_combout\ : std_logic;
SIGNAL \Mux113~9_combout\ : std_logic;
SIGNAL \Mux113~0_combout\ : std_logic;
SIGNAL \Mux113~26_combout\ : std_logic;
SIGNAL \RegFile[22][9]~q\ : std_logic;
SIGNAL \RegFile[17][9]~q\ : std_logic;
SIGNAL \Mux113~18_combout\ : std_logic;
SIGNAL \Mux113~5_combout\ : std_logic;
SIGNAL \Mux113~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[9]~12_combout\ : std_logic;
SIGNAL \Add2~33_OTERM719_OTERM823\ : std_logic;
SIGNAL \Add1~38\ : std_logic;
SIGNAL \Add1~42\ : std_logic;
SIGNAL \Add1~46\ : std_logic;
SIGNAL \Add1~50\ : std_logic;
SIGNAL \Add1~54\ : std_logic;
SIGNAL \Add1~57_sumout\ : std_logic;
SIGNAL \avm_d_readdata[22]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[14]~1_RESYN1094_BDD1095\ : std_logic;
SIGNAL \Comb:vRegWriteData[14]~1_RESYN1096_BDD1097\ : std_logic;
SIGNAL \Comb:vRegWriteData[14]~1_combout\ : std_logic;
SIGNAL \RegFile[29][14]~q\ : std_logic;
SIGNAL \RegFile[30][14]~feeder_combout\ : std_logic;
SIGNAL \RegFile[30][14]~q\ : std_logic;
SIGNAL \RegFile[31][14]~q\ : std_logic;
SIGNAL \RegFile[25][14]~q\ : std_logic;
SIGNAL \RegFile[27][14]~feeder_combout\ : std_logic;
SIGNAL \RegFile[27][14]~q\ : std_logic;
SIGNAL \RegFile[26][14]~feeder_combout\ : std_logic;
SIGNAL \RegFile[26][14]~q\ : std_logic;
SIGNAL \RegFile[24][14]~feeder_combout\ : std_logic;
SIGNAL \RegFile[24][14]~q\ : std_logic;
SIGNAL \Mux108~22_combout\ : std_logic;
SIGNAL \RegFile[28][14]~q\ : std_logic;
SIGNAL \Mux108~9_combout\ : std_logic;
SIGNAL \RegFile[21][14]~feeder_combout\ : std_logic;
SIGNAL \RegFile[21][14]~q\ : std_logic;
SIGNAL \RegFile[22][14]~q\ : std_logic;
SIGNAL \RegFile[23][14]~q\ : std_logic;
SIGNAL \RegFile[17][14]~q\ : std_logic;
SIGNAL \RegFile[19][14]~q\ : std_logic;
SIGNAL \RegFile[18][14]~q\ : std_logic;
SIGNAL \RegFile[16][14]~q\ : std_logic;
SIGNAL \Mux108~18_combout\ : std_logic;
SIGNAL \RegFile[20][14]~feeder_combout\ : std_logic;
SIGNAL \RegFile[20][14]~q\ : std_logic;
SIGNAL \Mux108~5_combout\ : std_logic;
SIGNAL \RegFile[3][14]~q\ : std_logic;
SIGNAL \RegFile[2][14]~q\ : std_logic;
SIGNAL \RegFile[7][14]~q\ : std_logic;
SIGNAL \RegFile[5][14]~feeder_combout\ : std_logic;
SIGNAL \RegFile[5][14]~q\ : std_logic;
SIGNAL \RegFile[4][14]~feeder_combout\ : std_logic;
SIGNAL \RegFile[4][14]~q\ : std_logic;
SIGNAL \RegFile[6][14]~q\ : std_logic;
SIGNAL \Mux108~0_combout\ : std_logic;
SIGNAL \RegFile[1][14]~feeder_combout\ : std_logic;
SIGNAL \RegFile[1][14]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux108~26_combout\ : std_logic;
SIGNAL \RegFile[15][14]~q\ : std_logic;
SIGNAL \RegFile[13][14]~q\ : std_logic;
SIGNAL \RegFile[14][14]~feeder_combout\ : std_logic;
SIGNAL \RegFile[14][14]~q\ : std_logic;
SIGNAL \RegFile[9][14]~q\ : std_logic;
SIGNAL \RegFile[10][14]~feeder_combout\ : std_logic;
SIGNAL \RegFile[10][14]~q\ : std_logic;
SIGNAL \RegFile[11][14]~q\ : std_logic;
SIGNAL \RegFile[8][14]~feeder_combout\ : std_logic;
SIGNAL \RegFile[8][14]~q\ : std_logic;
SIGNAL \Mux108~14_combout\ : std_logic;
SIGNAL \RegFile[12][14]~feeder_combout\ : std_logic;
SIGNAL \RegFile[12][14]~q\ : std_logic;
SIGNAL \Mux108~1_combout\ : std_logic;
SIGNAL \Mux108~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[14]~7_combout\ : std_logic;
SIGNAL \Add2~57_OTERM707_OTERM815\ : std_logic;
SIGNAL \Add2~58\ : std_logic;
SIGNAL \Add2~61_sumout\ : std_logic;
SIGNAL \ShiftRight1~54_combout\ : std_logic;
SIGNAL \Selector17~1_combout\ : std_logic;
SIGNAL \Selector17~2_combout\ : std_logic;
SIGNAL \Selector17~3_combout\ : std_logic;
SIGNAL \Selector17~5_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[15]~1_RESYN1048_BDD1049\ : std_logic;
SIGNAL \Comb:vRegWriteData[15]~1_RESYN1046_BDD1047\ : std_logic;
SIGNAL \Comb:vRegWriteData[15]~1_combout\ : std_logic;
SIGNAL \RegFile[31][15]~q\ : std_logic;
SIGNAL \Mux107~22_combout\ : std_logic;
SIGNAL \Mux107~9_combout\ : std_logic;
SIGNAL \Mux107~14_combout\ : std_logic;
SIGNAL \Mux107~1_combout\ : std_logic;
SIGNAL \Mux107~18_combout\ : std_logic;
SIGNAL \Mux107~5_combout\ : std_logic;
SIGNAL \RegFile[6][15]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux107~0_combout\ : std_logic;
SIGNAL \Mux107~26_combout\ : std_logic;
SIGNAL \Mux107~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[15]~6_combout\ : std_logic;
SIGNAL \Add1~61_sumout\ : std_logic;
SIGNAL \vAluRes~52_combout\ : std_logic;
SIGNAL \Add3~2\ : std_logic;
SIGNAL \Add3~6\ : std_logic;
SIGNAL \Add3~10\ : std_logic;
SIGNAL \Add3~14\ : std_logic;
SIGNAL \Add3~18\ : std_logic;
SIGNAL \Add3~22\ : std_logic;
SIGNAL \Add3~26\ : std_logic;
SIGNAL \Add3~30\ : std_logic;
SIGNAL \Add3~34\ : std_logic;
SIGNAL \Add3~38\ : std_logic;
SIGNAL \Add3~42\ : std_logic;
SIGNAL \Add3~46\ : std_logic;
SIGNAL \Add3~50\ : std_logic;
SIGNAL \Add3~54\ : std_logic;
SIGNAL \Add3~58\ : std_logic;
SIGNAL \Add3~61_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[15]~0_combout\ : std_logic;
SIGNAL \Mux44~0_combout\ : std_logic;
SIGNAL \NxR~10_combout\ : std_logic;
SIGNAL \NxR~9_combout\ : std_logic;
SIGNAL \NxR~11_combout\ : std_logic;
SIGNAL \R.incPC~q\ : std_logic;
SIGNAL \NxR.curPC[31]~0_combout\ : std_logic;
SIGNAL \Add0~54\ : std_logic;
SIGNAL \Add0~58\ : std_logic;
SIGNAL \Add0~61_sumout\ : std_logic;
SIGNAL \R.regWriteData[17]~feeder_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[17]~1_RESYN1124_BDD1125\ : std_logic;
SIGNAL \avm_d_readdata[9]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[17]~1_RESYN1120_BDD1121\ : std_logic;
SIGNAL \Comb:vRegWriteData[17]~1_RESYN1122_BDD1123\ : std_logic;
SIGNAL \Comb:vRegWriteData[17]~1_combout\ : std_logic;
SIGNAL \RegFile[13][17]~q\ : std_logic;
SIGNAL \Mux105~14_combout\ : std_logic;
SIGNAL \Mux105~1_combout\ : std_logic;
SIGNAL \Mux105~18_combout\ : std_logic;
SIGNAL \Mux105~5_combout\ : std_logic;
SIGNAL \Mux105~0_combout\ : std_logic;
SIGNAL \RegFile[1][17]~q\ : std_logic;
SIGNAL \Mux105~26_combout\ : std_logic;
SIGNAL \Mux105~22_combout\ : std_logic;
SIGNAL \Mux105~9_combout\ : std_logic;
SIGNAL \Mux105~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[17]~4_combout\ : std_logic;
SIGNAL \Add2~65_OTERM703_OTERM807\ : std_logic;
SIGNAL \Add2~69_sumout\ : std_logic;
SIGNAL \Selector15~5_combout\ : std_logic;
SIGNAL \Add3~62\ : std_logic;
SIGNAL \Add3~66\ : std_logic;
SIGNAL \Add3~69_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[17]~0_combout\ : std_logic;
SIGNAL \Add0~62\ : std_logic;
SIGNAL \Add0~65_sumout\ : std_logic;
SIGNAL \R.regWriteData[18]~feeder_combout\ : std_logic;
SIGNAL \Add1~73_sumout\ : std_logic;
SIGNAL \Add2~73_sumout\ : std_logic;
SIGNAL \avm_d_readdata[10]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[18]~1_RESYN1736_BDD1737\ : std_logic;
SIGNAL \Comb:vRegWriteData[18]~1_RESYN1738_BDD1739\ : std_logic;
SIGNAL \Comb:vRegWriteData[18]~1_RESYN1740_BDD1741\ : std_logic;
SIGNAL \Comb:vRegWriteData[18]~1_combout\ : std_logic;
SIGNAL \RegFile[21][18]~q\ : std_logic;
SIGNAL \Mux72~18_combout\ : std_logic;
SIGNAL \Mux72~5_combout\ : std_logic;
SIGNAL \RegFile[4][18]~q\ : std_logic;
SIGNAL \RegFile[6][18]~q\ : std_logic;
SIGNAL \Mux72~0_combout\ : std_logic;
SIGNAL \Mux72~26_combout\ : std_logic;
SIGNAL \RegFile[30][18]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux72~22_combout\ : std_logic;
SIGNAL \Mux72~9_combout\ : std_logic;
SIGNAL \RegFile[10][18]~q\ : std_logic;
SIGNAL \Mux72~14_combout\ : std_logic;
SIGNAL \Mux72~1_combout\ : std_logic;
SIGNAL \Mux72~13_combout\ : std_logic;
SIGNAL \Mux236~0_combout\ : std_logic;
SIGNAL \Selector14~1_combout\ : std_logic;
SIGNAL \Selector14~2_combout\ : std_logic;
SIGNAL \Selector14~3_combout\ : std_logic;
SIGNAL \Add3~70\ : std_logic;
SIGNAL \Add3~73_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[18]~0_combout\ : std_logic;
SIGNAL \Add0~66\ : std_logic;
SIGNAL \Add0~69_sumout\ : std_logic;
SIGNAL \R.regWriteData[19]~feeder_combout\ : std_logic;
SIGNAL \avm_d_readdata[11]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[19]~0_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[19]~1_combout\ : std_logic;
SIGNAL \RegFile[3][19]~q\ : std_logic;
SIGNAL \Mux71~0_combout\ : std_logic;
SIGNAL \RegFile[1][19]~q\ : std_logic;
SIGNAL \Mux71~26_combout\ : std_logic;
SIGNAL \Mux71~22_combout\ : std_logic;
SIGNAL \Mux71~9_combout\ : std_logic;
SIGNAL \Mux71~14_combout\ : std_logic;
SIGNAL \Mux71~1_combout\ : std_logic;
SIGNAL \Mux71~18_combout\ : std_logic;
SIGNAL \Mux71~5_combout\ : std_logic;
SIGNAL \Mux71~13_combout\ : std_logic;
SIGNAL \Mux235~0_combout\ : std_logic;
SIGNAL \Add2~78\ : std_logic;
SIGNAL \Add2~81_sumout\ : std_logic;
SIGNAL \avm_d_readdata[12]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[20]~1_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[20]~2_RESYN1110_BDD1111\ : std_logic;
SIGNAL \Comb:vRegWriteData[20]~2_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[20]~0_combout\ : std_logic;
SIGNAL \RegFile[6][20]~q\ : std_logic;
SIGNAL \RegFile[7][20]~q\ : std_logic;
SIGNAL \RegFile[4][20]~q\ : std_logic;
SIGNAL \RegFile[5][20]~feeder_combout\ : std_logic;
SIGNAL \RegFile[5][20]~q\ : std_logic;
SIGNAL \Mux102~0_combout\ : std_logic;
SIGNAL \RegFile[3][20]~q\ : std_logic;
SIGNAL \RegFile[2][20]~q\ : std_logic;
SIGNAL \RegFile[1][20]~feeder_combout\ : std_logic;
SIGNAL \RegFile[1][20]~q\ : std_logic;
SIGNAL \Mux102~26_combout\ : std_logic;
SIGNAL \RegFile[21][20]~q\ : std_logic;
SIGNAL \RegFile[23][20]~q\ : std_logic;
SIGNAL \RegFile[22][20]~q\ : std_logic;
SIGNAL \RegFile[17][20]~q\ : std_logic;
SIGNAL \RegFile[18][20]~feeder_combout\ : std_logic;
SIGNAL \RegFile[18][20]~q\ : std_logic;
SIGNAL \RegFile[19][20]~q\ : std_logic;
SIGNAL \RegFile[16][20]~feeder_combout\ : std_logic;
SIGNAL \RegFile[16][20]~q\ : std_logic;
SIGNAL \Mux102~18_combout\ : std_logic;
SIGNAL \RegFile[20][20]~q\ : std_logic;
SIGNAL \Mux102~5_combout\ : std_logic;
SIGNAL \RegFile[15][20]~q\ : std_logic;
SIGNAL \RegFile[13][20]~q\ : std_logic;
SIGNAL \RegFile[14][20]~DUPLICATE_q\ : std_logic;
SIGNAL \RegFile[11][20]~q\ : std_logic;
SIGNAL \RegFile[10][20]~feeder_combout\ : std_logic;
SIGNAL \RegFile[10][20]~q\ : std_logic;
SIGNAL \RegFile[9][20]~q\ : std_logic;
SIGNAL \RegFile[8][20]~feeder_combout\ : std_logic;
SIGNAL \RegFile[8][20]~q\ : std_logic;
SIGNAL \Mux102~14_combout\ : std_logic;
SIGNAL \RegFile[12][20]~q\ : std_logic;
SIGNAL \Mux102~1_combout\ : std_logic;
SIGNAL \RegFile[31][20]~q\ : std_logic;
SIGNAL \RegFile[29][20]~q\ : std_logic;
SIGNAL \RegFile[30][20]~feeder_combout\ : std_logic;
SIGNAL \RegFile[30][20]~q\ : std_logic;
SIGNAL \RegFile[25][20]~q\ : std_logic;
SIGNAL \RegFile[26][20]~feeder_combout\ : std_logic;
SIGNAL \RegFile[26][20]~q\ : std_logic;
SIGNAL \RegFile[27][20]~q\ : std_logic;
SIGNAL \RegFile[24][20]~feeder_combout\ : std_logic;
SIGNAL \RegFile[24][20]~q\ : std_logic;
SIGNAL \Mux102~22_combout\ : std_logic;
SIGNAL \RegFile[28][20]~feeder_combout\ : std_logic;
SIGNAL \RegFile[28][20]~q\ : std_logic;
SIGNAL \Mux102~9_combout\ : std_logic;
SIGNAL \Mux102~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[20]~1_combout\ : std_logic;
SIGNAL \Add2~82\ : std_logic;
SIGNAL \Add2~86\ : std_logic;
SIGNAL \Add2~90\ : std_logic;
SIGNAL \Add2~94\ : std_logic;
SIGNAL \Add2~98\ : std_logic;
SIGNAL \Add2~102\ : std_logic;
SIGNAL \Add2~106\ : std_logic;
SIGNAL \Add2~110\ : std_logic;
SIGNAL \Add2~114\ : std_logic;
SIGNAL \Add2~118\ : std_logic;
SIGNAL \Add2~121_sumout\ : std_logic;
SIGNAL \Selector2~3_combout\ : std_logic;
SIGNAL \avm_d_readdata[6]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[30]~1_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[30]~2_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[30]~0_combout\ : std_logic;
SIGNAL \RegFile[23][30]~q\ : std_logic;
SIGNAL \Mux60~18_combout\ : std_logic;
SIGNAL \Mux60~5_combout\ : std_logic;
SIGNAL \RegFile[30][30]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux60~22_combout\ : std_logic;
SIGNAL \Mux60~9_combout\ : std_logic;
SIGNAL \Mux60~0_combout\ : std_logic;
SIGNAL \Mux60~26_combout\ : std_logic;
SIGNAL \Mux60~14_combout\ : std_logic;
SIGNAL \Mux60~1_combout\ : std_logic;
SIGNAL \Mux60~13_combout\ : std_logic;
SIGNAL \Mux224~0_combout\ : std_logic;
SIGNAL \ShiftRight0~0_combout\ : std_logic;
SIGNAL \ShiftRight0~0_OTERM17\ : std_logic;
SIGNAL \Selector7~0_combout\ : std_logic;
SIGNAL \ShiftLeft0~42_combout\ : std_logic;
SIGNAL \ShiftLeft0~42_OTERM41\ : std_logic;
SIGNAL \ShiftLeft0~43_combout\ : std_logic;
SIGNAL \Selector7~1_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[25]~3_combout\ : std_logic;
SIGNAL \avm_d_readdata[1]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[25]~1_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[25]~2_RESYN1106_BDD1107\ : std_logic;
SIGNAL \Comb:vRegWriteData[25]~2_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[25]~0_combout\ : std_logic;
SIGNAL \RegFile[31][25]~q\ : std_logic;
SIGNAL \Mux65~22_combout\ : std_logic;
SIGNAL \Mux65~9_combout\ : std_logic;
SIGNAL \Mux65~18_combout\ : std_logic;
SIGNAL \Mux65~5_combout\ : std_logic;
SIGNAL \Mux65~0_combout\ : std_logic;
SIGNAL \Mux65~26_combout\ : std_logic;
SIGNAL \Mux65~14_combout\ : std_logic;
SIGNAL \Mux65~1_combout\ : std_logic;
SIGNAL \Mux65~13_combout\ : std_logic;
SIGNAL \Mux229~0_combout\ : std_logic;
SIGNAL \Add1~102\ : std_logic;
SIGNAL \Add1~106\ : std_logic;
SIGNAL \Add1~110\ : std_logic;
SIGNAL \Add1~114\ : std_logic;
SIGNAL \Add1~117_sumout\ : std_logic;
SIGNAL \Selector3~3_combout\ : std_logic;
SIGNAL \avm_d_readdata[5]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[29]~1_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[29]~2_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[29]~0_combout\ : std_logic;
SIGNAL \RegFile[31][29]~q\ : std_logic;
SIGNAL \RegFile[30][29]~feeder_combout\ : std_logic;
SIGNAL \RegFile[30][29]~q\ : std_logic;
SIGNAL \RegFile[29][29]~q\ : std_logic;
SIGNAL \RegFile[27][29]~q\ : std_logic;
SIGNAL \RegFile[25][29]~q\ : std_logic;
SIGNAL \RegFile[26][29]~q\ : std_logic;
SIGNAL \RegFile[24][29]~feeder_combout\ : std_logic;
SIGNAL \RegFile[24][29]~q\ : std_logic;
SIGNAL \Mux93~22_combout\ : std_logic;
SIGNAL \RegFile[28][29]~feeder_combout\ : std_logic;
SIGNAL \RegFile[28][29]~q\ : std_logic;
SIGNAL \Mux93~9_combout\ : std_logic;
SIGNAL \RegFile[23][29]~q\ : std_logic;
SIGNAL \RegFile[22][29]~feeder_combout\ : std_logic;
SIGNAL \RegFile[22][29]~q\ : std_logic;
SIGNAL \RegFile[21][29]~q\ : std_logic;
SIGNAL \RegFile[19][29]~q\ : std_logic;
SIGNAL \RegFile[17][29]~q\ : std_logic;
SIGNAL \RegFile[18][29]~feeder_combout\ : std_logic;
SIGNAL \RegFile[18][29]~q\ : std_logic;
SIGNAL \RegFile[16][29]~q\ : std_logic;
SIGNAL \Mux93~18_combout\ : std_logic;
SIGNAL \RegFile[20][29]~feeder_combout\ : std_logic;
SIGNAL \RegFile[20][29]~q\ : std_logic;
SIGNAL \Mux93~5_combout\ : std_logic;
SIGNAL \RegFile[3][29]~q\ : std_logic;
SIGNAL \RegFile[2][29]~q\ : std_logic;
SIGNAL \RegFile[7][29]~q\ : std_logic;
SIGNAL \RegFile[4][29]~feeder_combout\ : std_logic;
SIGNAL \RegFile[4][29]~q\ : std_logic;
SIGNAL \RegFile[6][29]~q\ : std_logic;
SIGNAL \RegFile[5][29]~q\ : std_logic;
SIGNAL \Mux93~0_combout\ : std_logic;
SIGNAL \RegFile[1][29]~q\ : std_logic;
SIGNAL \Mux93~26_combout\ : std_logic;
SIGNAL \RegFile[13][29]~feeder_combout\ : std_logic;
SIGNAL \RegFile[13][29]~q\ : std_logic;
SIGNAL \RegFile[14][29]~feeder_combout\ : std_logic;
SIGNAL \RegFile[14][29]~q\ : std_logic;
SIGNAL \RegFile[15][29]~q\ : std_logic;
SIGNAL \RegFile[11][29]~q\ : std_logic;
SIGNAL \RegFile[10][29]~feeder_combout\ : std_logic;
SIGNAL \RegFile[10][29]~q\ : std_logic;
SIGNAL \RegFile[9][29]~q\ : std_logic;
SIGNAL \RegFile[8][29]~q\ : std_logic;
SIGNAL \Mux93~14_combout\ : std_logic;
SIGNAL \RegFile[12][29]~q\ : std_logic;
SIGNAL \Mux93~1_combout\ : std_logic;
SIGNAL \Mux93~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[29]~31_combout\ : std_logic;
SIGNAL \Selector3~1_combout\ : std_logic;
SIGNAL \ShiftLeft0~19_combout\ : std_logic;
SIGNAL \ShiftLeft0~51_combout\ : std_logic;
SIGNAL \ShiftLeft0~51_OTERM763\ : std_logic;
SIGNAL \ShiftLeft0~52_combout\ : std_logic;
SIGNAL \Selector3~0_combout\ : std_logic;
SIGNAL \Selector3~2_combout\ : std_logic;
SIGNAL \Comb:vJumpAdr[29]~0_RESYN1034_BDD1035\ : std_logic;
SIGNAL \Mux126~0_combout\ : std_logic;
SIGNAL \Mux133~0_combout\ : std_logic;
SIGNAL \Add3~74\ : std_logic;
SIGNAL \Add3~78\ : std_logic;
SIGNAL \Add3~82\ : std_logic;
SIGNAL \Add3~86\ : std_logic;
SIGNAL \Add3~90\ : std_logic;
SIGNAL \Add3~94\ : std_logic;
SIGNAL \Add3~98\ : std_logic;
SIGNAL \Add3~102\ : std_logic;
SIGNAL \Add3~106\ : std_logic;
SIGNAL \Add3~110\ : std_logic;
SIGNAL \Add3~114\ : std_logic;
SIGNAL \Add3~117_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[29]~0_combout\ : std_logic;
SIGNAL \Mux61~22_combout\ : std_logic;
SIGNAL \Mux61~9_combout\ : std_logic;
SIGNAL \Mux61~18_combout\ : std_logic;
SIGNAL \Mux61~5_combout\ : std_logic;
SIGNAL \Mux61~14_combout\ : std_logic;
SIGNAL \Mux61~1_combout\ : std_logic;
SIGNAL \Mux61~0_combout\ : std_logic;
SIGNAL \RegFile[1][29]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux61~26_combout\ : std_logic;
SIGNAL \Mux61~13_combout\ : std_logic;
SIGNAL \Mux225~0_combout\ : std_logic;
SIGNAL \ShiftRight1~13_combout\ : std_logic;
SIGNAL \ShiftRight1~13_OTERM15\ : std_logic;
SIGNAL \ShiftRight1~41_combout\ : std_logic;
SIGNAL \Selector27~5_combout\ : std_logic;
SIGNAL \vAluRes~5_RESYN1070_BDD1071\ : std_logic;
SIGNAL \vAluRes~5_combout\ : std_logic;
SIGNAL \Add3~21_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[5]~0_combout\ : std_logic;
SIGNAL \Add0~14\ : std_logic;
SIGNAL \Add0~18\ : std_logic;
SIGNAL \Add0~21_sumout\ : std_logic;
SIGNAL \R.regWriteData[7]~feeder_combout\ : std_logic;
SIGNAL \vAluRes~7_RESYN1076_RESYN1132_BDD1133\ : std_logic;
SIGNAL \vAluRes~7_RESYN1076_BDD1077\ : std_logic;
SIGNAL \Comb:vRegWriteData[7]~0_RESYN1118_BDD1119\ : std_logic;
SIGNAL \Comb:vRegWriteData[7]~0_combout\ : std_logic;
SIGNAL \RegFile[2][7]~feeder_combout\ : std_logic;
SIGNAL \RegFile[2][7]~q\ : std_logic;
SIGNAL \Mux115~0_combout\ : std_logic;
SIGNAL \Mux115~26_combout\ : std_logic;
SIGNAL \Mux115~18_combout\ : std_logic;
SIGNAL \Mux115~5_combout\ : std_logic;
SIGNAL \Mux115~14_combout\ : std_logic;
SIGNAL \Mux115~1_combout\ : std_logic;
SIGNAL \RegFile[30][7]~q\ : std_logic;
SIGNAL \Mux115~22_combout\ : std_logic;
SIGNAL \Mux115~9_combout\ : std_logic;
SIGNAL \Mux115~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[7]~14_combout\ : std_logic;
SIGNAL \Add2~25_OTERM723_OTERM831\ : std_logic;
SIGNAL \Add1~29_sumout\ : std_logic;
SIGNAL \vAluRes~7_combout\ : std_logic;
SIGNAL \Add3~29_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[7]~0_combout\ : std_logic;
SIGNAL \Add0~22\ : std_logic;
SIGNAL \Add0~25_sumout\ : std_logic;
SIGNAL \R.regWriteData[8]~feeder_combout\ : std_logic;
SIGNAL \Selector24~0_RTM0421_combout\ : std_logic;
SIGNAL \Selector24~0_OTERM419\ : std_logic;
SIGNAL \Selector24~1_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[8]~1_RESYN1734_BDD1735\ : std_logic;
SIGNAL \ShiftLeft0~11_combout\ : std_logic;
SIGNAL \ShiftRight0~10_combout\ : std_logic;
SIGNAL \ShiftRight1~7_combout\ : std_logic;
SIGNAL \ShiftRight1~7_OTERM259\ : std_logic;
SIGNAL \ShiftRight1~46_combout\ : std_logic;
SIGNAL \Selector24~3_combout\ : std_logic;
SIGNAL \Add2~33_sumout\ : std_logic;
SIGNAL \avm_d_readdata[16]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[8]~1_RESYN1730_BDD1731\ : std_logic;
SIGNAL \Comb:vRegWriteData[8]~1_RESYN1732_BDD1733\ : std_logic;
SIGNAL \Comb:vRegWriteData[8]~1_combout\ : std_logic;
SIGNAL \RegFile[3][8]~q\ : std_logic;
SIGNAL \RegFile[2][8]~q\ : std_logic;
SIGNAL \RegFile[5][8]~feeder_combout\ : std_logic;
SIGNAL \RegFile[5][8]~q\ : std_logic;
SIGNAL \RegFile[6][8]~feeder_combout\ : std_logic;
SIGNAL \RegFile[6][8]~DUPLICATE_q\ : std_logic;
SIGNAL \RegFile[4][8]~q\ : std_logic;
SIGNAL \RegFile[7][8]~q\ : std_logic;
SIGNAL \Mux114~0_combout\ : std_logic;
SIGNAL \RegFile[1][8]~feeder_combout\ : std_logic;
SIGNAL \RegFile[1][8]~q\ : std_logic;
SIGNAL \Mux114~26_combout\ : std_logic;
SIGNAL \RegFile[13][8]~q\ : std_logic;
SIGNAL \RegFile[14][8]~q\ : std_logic;
SIGNAL \RegFile[15][8]~q\ : std_logic;
SIGNAL \RegFile[9][8]~q\ : std_logic;
SIGNAL \RegFile[11][8]~feeder_combout\ : std_logic;
SIGNAL \RegFile[11][8]~DUPLICATE_q\ : std_logic;
SIGNAL \RegFile[10][8]~feeder_combout\ : std_logic;
SIGNAL \RegFile[10][8]~q\ : std_logic;
SIGNAL \RegFile[8][8]~feeder_combout\ : std_logic;
SIGNAL \RegFile[8][8]~q\ : std_logic;
SIGNAL \Mux114~14_combout\ : std_logic;
SIGNAL \RegFile[12][8]~feeder_combout\ : std_logic;
SIGNAL \RegFile[12][8]~q\ : std_logic;
SIGNAL \Mux114~1_combout\ : std_logic;
SIGNAL \RegFile[21][8]~q\ : std_logic;
SIGNAL \RegFile[23][8]~q\ : std_logic;
SIGNAL \RegFile[22][8]~feeder_combout\ : std_logic;
SIGNAL \RegFile[22][8]~q\ : std_logic;
SIGNAL \RegFile[17][8]~q\ : std_logic;
SIGNAL \RegFile[19][8]~q\ : std_logic;
SIGNAL \RegFile[18][8]~feeder_combout\ : std_logic;
SIGNAL \RegFile[18][8]~q\ : std_logic;
SIGNAL \RegFile[16][8]~feeder_combout\ : std_logic;
SIGNAL \RegFile[16][8]~q\ : std_logic;
SIGNAL \Mux114~18_combout\ : std_logic;
SIGNAL \RegFile[20][8]~feeder_combout\ : std_logic;
SIGNAL \RegFile[20][8]~q\ : std_logic;
SIGNAL \Mux114~5_combout\ : std_logic;
SIGNAL \RegFile[29][8]~q\ : std_logic;
SIGNAL \RegFile[31][8]~feeder_combout\ : std_logic;
SIGNAL \RegFile[31][8]~DUPLICATE_q\ : std_logic;
SIGNAL \RegFile[30][8]~feeder_combout\ : std_logic;
SIGNAL \RegFile[30][8]~q\ : std_logic;
SIGNAL \RegFile[27][8]~q\ : std_logic;
SIGNAL \RegFile[26][8]~q\ : std_logic;
SIGNAL \RegFile[25][8]~feeder_combout\ : std_logic;
SIGNAL \RegFile[25][8]~q\ : std_logic;
SIGNAL \RegFile[24][8]~feeder_combout\ : std_logic;
SIGNAL \RegFile[24][8]~q\ : std_logic;
SIGNAL \Mux114~22_combout\ : std_logic;
SIGNAL \RegFile[28][8]~feeder_combout\ : std_logic;
SIGNAL \RegFile[28][8]~q\ : std_logic;
SIGNAL \Mux114~9_combout\ : std_logic;
SIGNAL \Mux114~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[8]~13_combout\ : std_logic;
SIGNAL \Add2~33_OTERM719_OTERM827\ : std_logic;
SIGNAL \Add1~33_sumout\ : std_logic;
SIGNAL \Selector24~4_combout\ : std_logic;
SIGNAL \vAluRes~31_combout\ : std_logic;
SIGNAL \vAluRes~8_combout\ : std_logic;
SIGNAL \Add3~33_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[8]~0_combout\ : std_logic;
SIGNAL \RegFile[31][8]~q\ : std_logic;
SIGNAL \Mux82~22_combout\ : std_logic;
SIGNAL \Mux82~9_combout\ : std_logic;
SIGNAL \RegFile[6][8]~q\ : std_logic;
SIGNAL \Mux82~0_combout\ : std_logic;
SIGNAL \Mux82~26_combout\ : std_logic;
SIGNAL \RegFile[11][8]~q\ : std_logic;
SIGNAL \Mux82~14_combout\ : std_logic;
SIGNAL \Mux82~1_combout\ : std_logic;
SIGNAL \RegFile[18][8]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux82~18_combout\ : std_logic;
SIGNAL \Mux82~5_combout\ : std_logic;
SIGNAL \Mux82~13_combout\ : std_logic;
SIGNAL \Mux246~0_combout\ : std_logic;
SIGNAL \ShiftLeft0~14_combout\ : std_logic;
SIGNAL \ShiftLeft0~14_OTERM753\ : std_logic;
SIGNAL \ShiftLeft0~31_combout\ : std_logic;
SIGNAL \ShiftRight1~33_combout\ : std_logic;
SIGNAL \ShiftRight0~5_combout\ : std_logic;
SIGNAL \Selector13~0_combout\ : std_logic;
SIGNAL \Selector13~2_combout\ : std_logic;
SIGNAL \Add3~77_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[19]~0_combout\ : std_logic;
SIGNAL \Add0~70\ : std_logic;
SIGNAL \Add0~74\ : std_logic;
SIGNAL \Add0~78\ : std_logic;
SIGNAL \Add0~82\ : std_logic;
SIGNAL \Add0~86\ : std_logic;
SIGNAL \Add0~89_sumout\ : std_logic;
SIGNAL \ShiftLeft0~41_combout\ : std_logic;
SIGNAL \Selector8~0_combout\ : std_logic;
SIGNAL \Selector8~1_combout\ : std_logic;
SIGNAL \Selector8~2_combout\ : std_logic;
SIGNAL \Selector8~3_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[24]~4_combout\ : std_logic;
SIGNAL \Add1~97_sumout\ : std_logic;
SIGNAL \Comb:vRegWriteData[24]~2_combout\ : std_logic;
SIGNAL \avm_d_readdata[0]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[24]~3_RESYN1104_BDD1105\ : std_logic;
SIGNAL \Comb:vRegWriteData[24]~3_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[24]~0_combout\ : std_logic;
SIGNAL \RegFile[29][24]~q\ : std_logic;
SIGNAL \RegFile[31][24]~q\ : std_logic;
SIGNAL \RegFile[30][24]~feeder_combout\ : std_logic;
SIGNAL \RegFile[30][24]~q\ : std_logic;
SIGNAL \RegFile[25][24]~feeder_combout\ : std_logic;
SIGNAL \RegFile[25][24]~q\ : std_logic;
SIGNAL \RegFile[27][24]~q\ : std_logic;
SIGNAL \RegFile[26][24]~q\ : std_logic;
SIGNAL \RegFile[24][24]~feeder_combout\ : std_logic;
SIGNAL \RegFile[24][24]~q\ : std_logic;
SIGNAL \Mux98~22_combout\ : std_logic;
SIGNAL \RegFile[28][24]~q\ : std_logic;
SIGNAL \Mux98~9_combout\ : std_logic;
SIGNAL \RegFile[3][24]~q\ : std_logic;
SIGNAL \RegFile[2][24]~feeder_combout\ : std_logic;
SIGNAL \RegFile[2][24]~q\ : std_logic;
SIGNAL \RegFile[5][24]~feeder_combout\ : std_logic;
SIGNAL \RegFile[5][24]~q\ : std_logic;
SIGNAL \RegFile[7][24]~q\ : std_logic;
SIGNAL \RegFile[6][24]~q\ : std_logic;
SIGNAL \RegFile[4][24]~feeder_combout\ : std_logic;
SIGNAL \RegFile[4][24]~q\ : std_logic;
SIGNAL \Mux98~0_combout\ : std_logic;
SIGNAL \RegFile[1][24]~q\ : std_logic;
SIGNAL \Mux98~26_combout\ : std_logic;
SIGNAL \RegFile[13][24]~q\ : std_logic;
SIGNAL \RegFile[15][24]~q\ : std_logic;
SIGNAL \RegFile[14][24]~q\ : std_logic;
SIGNAL \RegFile[9][24]~q\ : std_logic;
SIGNAL \RegFile[10][24]~q\ : std_logic;
SIGNAL \RegFile[11][24]~q\ : std_logic;
SIGNAL \RegFile[8][24]~feeder_combout\ : std_logic;
SIGNAL \RegFile[8][24]~q\ : std_logic;
SIGNAL \Mux98~14_combout\ : std_logic;
SIGNAL \RegFile[12][24]~feeder_combout\ : std_logic;
SIGNAL \RegFile[12][24]~q\ : std_logic;
SIGNAL \Mux98~1_combout\ : std_logic;
SIGNAL \RegFile[23][24]~q\ : std_logic;
SIGNAL \RegFile[21][24]~q\ : std_logic;
SIGNAL \RegFile[22][24]~q\ : std_logic;
SIGNAL \RegFile[17][24]~q\ : std_logic;
SIGNAL \RegFile[19][24]~feeder_combout\ : std_logic;
SIGNAL \RegFile[19][24]~q\ : std_logic;
SIGNAL \RegFile[18][24]~feeder_combout\ : std_logic;
SIGNAL \RegFile[18][24]~q\ : std_logic;
SIGNAL \RegFile[16][24]~q\ : std_logic;
SIGNAL \Mux98~18_combout\ : std_logic;
SIGNAL \RegFile[20][24]~feeder_combout\ : std_logic;
SIGNAL \RegFile[20][24]~q\ : std_logic;
SIGNAL \Mux98~5_combout\ : std_logic;
SIGNAL \Mux98~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[24]~26_combout\ : std_logic;
SIGNAL \Add2~97_sumout\ : std_logic;
SIGNAL \Selector8~4_combout\ : std_logic;
SIGNAL \Add3~97_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[24]~0_combout\ : std_logic;
SIGNAL \Mux66~14_combout\ : std_logic;
SIGNAL \Mux66~1_combout\ : std_logic;
SIGNAL \Mux66~22_combout\ : std_logic;
SIGNAL \Mux66~9_combout\ : std_logic;
SIGNAL \Mux66~18_combout\ : std_logic;
SIGNAL \Mux66~5_combout\ : std_logic;
SIGNAL \Mux66~0_combout\ : std_logic;
SIGNAL \Mux66~26_combout\ : std_logic;
SIGNAL \Mux66~13_combout\ : std_logic;
SIGNAL \Mux230~0_combout\ : std_logic;
SIGNAL \ShiftRight1~26_combout\ : std_logic;
SIGNAL \ShiftRight1~26_OTERM37\ : std_logic;
SIGNAL \ShiftRight1~28_combout\ : std_logic;
SIGNAL \ShiftRight1~28_OTERM23\ : std_logic;
SIGNAL \ShiftRight1~43_combout\ : std_logic;
SIGNAL \Selector26~4_combout\ : std_logic;
SIGNAL \vAluRes~6_RESYN1072_BDD1073\ : std_logic;
SIGNAL \vAluRes~6_combout\ : std_logic;
SIGNAL \Add3~25_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[6]~0_combout\ : std_logic;
SIGNAL \Mux84~0_combout\ : std_logic;
SIGNAL \Mux84~26_combout\ : std_logic;
SIGNAL \Mux84~22_combout\ : std_logic;
SIGNAL \Mux84~9_combout\ : std_logic;
SIGNAL \Mux84~18_combout\ : std_logic;
SIGNAL \Mux84~5_combout\ : std_logic;
SIGNAL \RegFile[14][6]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux84~14_combout\ : std_logic;
SIGNAL \Mux84~1_combout\ : std_logic;
SIGNAL \Mux84~13_combout\ : std_logic;
SIGNAL \Mux248~0_combout\ : std_logic;
SIGNAL \ShiftLeft0~10_combout\ : std_logic;
SIGNAL \ShiftLeft0~10_OTERM211\ : std_logic;
SIGNAL \ShiftLeft0~25_combout\ : std_logic;
SIGNAL \Selector16~1_RTM0795_combout\ : std_logic;
SIGNAL \Selector16~1_OTERM793\ : std_logic;
SIGNAL \Selector16~2_combout\ : std_logic;
SIGNAL \ShiftRight1~4_combout\ : std_logic;
SIGNAL \Selector16~3_combout\ : std_logic;
SIGNAL \Selector16~5_combout\ : std_logic;
SIGNAL \Add3~65_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[16]~0_combout\ : std_logic;
SIGNAL \RegFile[14][16]~q\ : std_logic;
SIGNAL \Mux74~14_combout\ : std_logic;
SIGNAL \RegFile[12][16]~q\ : std_logic;
SIGNAL \Mux74~1_combout\ : std_logic;
SIGNAL \Mux74~18_combout\ : std_logic;
SIGNAL \RegFile[20][16]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux74~5_combout\ : std_logic;
SIGNAL \RegFile[5][16]~q\ : std_logic;
SIGNAL \Mux74~0_combout\ : std_logic;
SIGNAL \Mux74~26_combout\ : std_logic;
SIGNAL \Mux74~22_combout\ : std_logic;
SIGNAL \Mux74~9_combout\ : std_logic;
SIGNAL \Mux74~13_combout\ : std_logic;
SIGNAL \Mux238~0_combout\ : std_logic;
SIGNAL \ShiftRight1~18_combout\ : std_logic;
SIGNAL \ShiftRight1~18_OTERM269\ : std_logic;
SIGNAL \ShiftRight1~47_combout\ : std_logic;
SIGNAL \Selector23~5_combout\ : std_logic;
SIGNAL \Selector23~0_combout\ : std_logic;
SIGNAL \Add3~37_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[9]~0_combout\ : std_logic;
SIGNAL \Add0~30\ : std_logic;
SIGNAL \Add0~33_sumout\ : std_logic;
SIGNAL \R.regWriteData[10]~feeder_combout\ : std_logic;
SIGNAL \ShiftRight1~49_combout\ : std_logic;
SIGNAL \Selector22~3_combout\ : std_logic;
SIGNAL \Add1~41_sumout\ : std_logic;
SIGNAL \Selector22~4_combout\ : std_logic;
SIGNAL \Add2~41_sumout\ : std_logic;
SIGNAL \Selector22~2_combout\ : std_logic;
SIGNAL \Selector22~5_combout\ : std_logic;
SIGNAL \avm_d_readdata[18]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[10]~0_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[10]~1_combout\ : std_logic;
SIGNAL \RegFile[2][10]~q\ : std_logic;
SIGNAL \Mux112~0_combout\ : std_logic;
SIGNAL \Mux112~26_combout\ : std_logic;
SIGNAL \Mux112~22_combout\ : std_logic;
SIGNAL \Mux112~9_combout\ : std_logic;
SIGNAL \Mux112~18_combout\ : std_logic;
SIGNAL \Mux112~5_combout\ : std_logic;
SIGNAL \RegFile[10][10]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux112~14_combout\ : std_logic;
SIGNAL \RegFile[12][10]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux112~1_combout\ : std_logic;
SIGNAL \Mux112~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[10]~9_combout\ : std_logic;
SIGNAL \Selector22~1_RTM0429_combout\ : std_logic;
SIGNAL \Selector22~1_OTERM427\ : std_logic;
SIGNAL \vAluRes~32_combout\ : std_logic;
SIGNAL \vAluRes~10_combout\ : std_logic;
SIGNAL \Add3~41_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[10]~0_combout\ : std_logic;
SIGNAL \Add0~34\ : std_logic;
SIGNAL \Add0~37_sumout\ : std_logic;
SIGNAL \R.regWriteData[11]~feeder_combout\ : std_logic;
SIGNAL \Selector21~0_combout\ : std_logic;
SIGNAL \Selector21~1_combout\ : std_logic;
SIGNAL \ShiftRight0~7_OTERM233\ : std_logic;
SIGNAL \Selector21~2_combout\ : std_logic;
SIGNAL \ShiftRight1~50_combout\ : std_logic;
SIGNAL \Selector21~3_combout\ : std_logic;
SIGNAL \Add2~45_sumout\ : std_logic;
SIGNAL \Selector21~5_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[11]~1_RESYN1040_BDD1041\ : std_logic;
SIGNAL \avm_d_readdata[19]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[11]~1_RESYN1038_BDD1039\ : std_logic;
SIGNAL \Comb:vRegWriteData[11]~1_combout\ : std_logic;
SIGNAL \RegFile[29][11]~q\ : std_logic;
SIGNAL \Mux79~22_combout\ : std_logic;
SIGNAL \Mux79~9_combout\ : std_logic;
SIGNAL \Mux79~0_combout\ : std_logic;
SIGNAL \Mux79~26_combout\ : std_logic;
SIGNAL \Mux79~18_combout\ : std_logic;
SIGNAL \Mux79~5_combout\ : std_logic;
SIGNAL \RegFile[11][11]~q\ : std_logic;
SIGNAL \Mux79~14_combout\ : std_logic;
SIGNAL \Mux79~1_combout\ : std_logic;
SIGNAL \Mux79~13_combout\ : std_logic;
SIGNAL \Mux243~0_combout\ : std_logic;
SIGNAL \Add1~45_sumout\ : std_logic;
SIGNAL \vAluRes~60_combout\ : std_logic;
SIGNAL \Add3~45_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[11]~0_combout\ : std_logic;
SIGNAL \Add0~38\ : std_logic;
SIGNAL \Add0~41_sumout\ : std_logic;
SIGNAL \R.regWriteData[12]~feeder_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[12]~1_RESYN1088_BDD1089\ : std_logic;
SIGNAL \avm_d_readdata[20]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[12]~1_RESYN1086_BDD1087\ : std_logic;
SIGNAL \Comb:vRegWriteData[12]~1_combout\ : std_logic;
SIGNAL \RegFile[13][12]~feeder_combout\ : std_logic;
SIGNAL \RegFile[13][12]~q\ : std_logic;
SIGNAL \Mux78~14_combout\ : std_logic;
SIGNAL \Mux78~1_combout\ : std_logic;
SIGNAL \Mux78~0_combout\ : std_logic;
SIGNAL \RegFile[2][12]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux78~26_combout\ : std_logic;
SIGNAL \Mux78~18_combout\ : std_logic;
SIGNAL \Mux78~5_combout\ : std_logic;
SIGNAL \Mux78~22_combout\ : std_logic;
SIGNAL \Mux78~9_combout\ : std_logic;
SIGNAL \Mux78~13_combout\ : std_logic;
SIGNAL \Mux242~0_combout\ : std_logic;
SIGNAL \Add2~49_sumout\ : std_logic;
SIGNAL \Selector20~4_combout\ : std_logic;
SIGNAL \Add3~49_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[12]~0_combout\ : std_logic;
SIGNAL \Add0~42\ : std_logic;
SIGNAL \Add0~45_sumout\ : std_logic;
SIGNAL \R.regWriteData[13]~feeder_combout\ : std_logic;
SIGNAL \Add2~53_sumout\ : std_logic;
SIGNAL \R.aluData2[13]~DUPLICATE_q\ : std_logic;
SIGNAL \Selector19~2_combout\ : std_logic;
SIGNAL \ShiftRight1~52_combout\ : std_logic;
SIGNAL \Selector19~0_combout\ : std_logic;
SIGNAL \Selector19~1_OTERM751_OTERM803\ : std_logic;
SIGNAL \Selector19~1_combout\ : std_logic;
SIGNAL \Selector19~3_combout\ : std_logic;
SIGNAL \Selector19~5_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[13]~1_RESYN1044_BDD1045\ : std_logic;
SIGNAL \avm_d_readdata[21]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[13]~1_RESYN1042_BDD1043\ : std_logic;
SIGNAL \Comb:vRegWriteData[13]~1_combout\ : std_logic;
SIGNAL \RegFile[29][13]~feeder_combout\ : std_logic;
SIGNAL \RegFile[29][13]~q\ : std_logic;
SIGNAL \RegFile[30][13]~q\ : std_logic;
SIGNAL \RegFile[31][13]~q\ : std_logic;
SIGNAL \RegFile[27][13]~q\ : std_logic;
SIGNAL \RegFile[25][13]~q\ : std_logic;
SIGNAL \RegFile[26][13]~q\ : std_logic;
SIGNAL \RegFile[24][13]~q\ : std_logic;
SIGNAL \Mux109~22_combout\ : std_logic;
SIGNAL \RegFile[28][13]~feeder_combout\ : std_logic;
SIGNAL \RegFile[28][13]~q\ : std_logic;
SIGNAL \Mux109~9_combout\ : std_logic;
SIGNAL \RegFile[13][13]~q\ : std_logic;
SIGNAL \RegFile[14][13]~q\ : std_logic;
SIGNAL \RegFile[15][13]~q\ : std_logic;
SIGNAL \RegFile[11][13]~q\ : std_logic;
SIGNAL \RegFile[10][13]~feeder_combout\ : std_logic;
SIGNAL \RegFile[10][13]~q\ : std_logic;
SIGNAL \RegFile[9][13]~q\ : std_logic;
SIGNAL \RegFile[8][13]~q\ : std_logic;
SIGNAL \Mux109~14_combout\ : std_logic;
SIGNAL \RegFile[12][13]~feeder_combout\ : std_logic;
SIGNAL \RegFile[12][13]~q\ : std_logic;
SIGNAL \Mux109~1_combout\ : std_logic;
SIGNAL \RegFile[3][13]~q\ : std_logic;
SIGNAL \RegFile[2][13]~q\ : std_logic;
SIGNAL \RegFile[4][13]~q\ : std_logic;
SIGNAL \RegFile[7][13]~q\ : std_logic;
SIGNAL \RegFile[6][13]~q\ : std_logic;
SIGNAL \RegFile[5][13]~q\ : std_logic;
SIGNAL \Mux109~0_combout\ : std_logic;
SIGNAL \RegFile[1][13]~q\ : std_logic;
SIGNAL \Mux109~26_combout\ : std_logic;
SIGNAL \RegFile[23][13]~q\ : std_logic;
SIGNAL \RegFile[22][13]~q\ : std_logic;
SIGNAL \RegFile[21][13]~q\ : std_logic;
SIGNAL \RegFile[17][13]~q\ : std_logic;
SIGNAL \RegFile[18][13]~feeder_combout\ : std_logic;
SIGNAL \RegFile[18][13]~q\ : std_logic;
SIGNAL \RegFile[19][13]~q\ : std_logic;
SIGNAL \RegFile[16][13]~feeder_combout\ : std_logic;
SIGNAL \RegFile[16][13]~q\ : std_logic;
SIGNAL \Mux109~18_combout\ : std_logic;
SIGNAL \RegFile[20][13]~q\ : std_logic;
SIGNAL \Mux109~5_combout\ : std_logic;
SIGNAL \Mux109~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[13]~10_combout\ : std_logic;
SIGNAL \Add1~53_sumout\ : std_logic;
SIGNAL \vAluRes~56_combout\ : std_logic;
SIGNAL \Add3~53_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[13]~0_combout\ : std_logic;
SIGNAL \Mux77~14_combout\ : std_logic;
SIGNAL \Mux77~1_combout\ : std_logic;
SIGNAL \Mux77~18_combout\ : std_logic;
SIGNAL \Mux77~5_combout\ : std_logic;
SIGNAL \Mux77~22_combout\ : std_logic;
SIGNAL \Mux77~9_combout\ : std_logic;
SIGNAL \Mux77~0_combout\ : std_logic;
SIGNAL \Mux77~26_combout\ : std_logic;
SIGNAL \Mux77~13_combout\ : std_logic;
SIGNAL \Mux241~0_combout\ : std_logic;
SIGNAL \ShiftRight1~36_combout\ : std_logic;
SIGNAL \ShiftRight1~36_OTERM281\ : std_logic;
SIGNAL \ShiftRight1~34_combout\ : std_logic;
SIGNAL \ShiftRight1~38_OTERM439_OTERM745\ : std_logic;
SIGNAL \ShiftRight1~38_combout\ : std_logic;
SIGNAL \Selector29~2_combout\ : std_logic;
SIGNAL \Add2~13_sumout\ : std_logic;
SIGNAL \Add1~13_sumout\ : std_logic;
SIGNAL \Selector29~3_combout\ : std_logic;
SIGNAL \Selector29~4_combout\ : std_logic;
SIGNAL \vAluRes~3_RESYN1066_BDD1067\ : std_logic;
SIGNAL \vAluRes~3_combout\ : std_logic;
SIGNAL \Add3~13_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[3]~0_combout\ : std_logic;
SIGNAL \Add0~5_sumout\ : std_logic;
SIGNAL \R.regWriteData[3]~feeder_combout\ : std_logic;
SIGNAL \avm_d_readdata[27]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[3]~0_RESYN1084_BDD1085\ : std_logic;
SIGNAL \Comb:vRegWriteData[3]~0_combout\ : std_logic;
SIGNAL \RegFile[13][3]~q\ : std_logic;
SIGNAL \Mux119~14_combout\ : std_logic;
SIGNAL \Mux119~1_combout\ : std_logic;
SIGNAL \Mux119~22_combout\ : std_logic;
SIGNAL \Mux119~9_combout\ : std_logic;
SIGNAL \Mux119~18_combout\ : std_logic;
SIGNAL \Mux119~5_combout\ : std_logic;
SIGNAL \Mux119~0_combout\ : std_logic;
SIGNAL \Mux119~26_combout\ : std_logic;
SIGNAL \Mux119~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[3]~18_combout\ : std_logic;
SIGNAL \Selector7~2_combout\ : std_logic;
SIGNAL \Selector7~5_combout\ : std_logic;
SIGNAL \Selector7~4_combout\ : std_logic;
SIGNAL \vAluRes~25_combout\ : std_logic;
SIGNAL \Add3~101_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[25]~0_combout\ : std_logic;
SIGNAL \Add0~94\ : std_logic;
SIGNAL \Add0~97_sumout\ : std_logic;
SIGNAL \avm_d_readdata[2]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[26]~1_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[26]~2_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[26]~0_combout\ : std_logic;
SIGNAL \RegFile[21][26]~q\ : std_logic;
SIGNAL \Mux64~18_combout\ : std_logic;
SIGNAL \Mux64~5_combout\ : std_logic;
SIGNAL \RegFile[2][26]~DUPLICATE_q\ : std_logic;
SIGNAL \RegFile[7][26]~q\ : std_logic;
SIGNAL \Mux64~0_combout\ : std_logic;
SIGNAL \Mux64~26_combout\ : std_logic;
SIGNAL \Mux64~22_combout\ : std_logic;
SIGNAL \Mux64~9_combout\ : std_logic;
SIGNAL \RegFile[10][26]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux64~14_combout\ : std_logic;
SIGNAL \Mux64~1_combout\ : std_logic;
SIGNAL \Mux64~13_combout\ : std_logic;
SIGNAL \Mux228~0_combout\ : std_logic;
SIGNAL \ShiftRight1~12_combout\ : std_logic;
SIGNAL \ShiftRight1~12_OTERM57\ : std_logic;
SIGNAL \ShiftRight0~1_combout\ : std_logic;
SIGNAL \ShiftRight1~15_combout\ : std_logic;
SIGNAL \ShiftRight1~15_OTERM199\ : std_logic;
SIGNAL \ShiftRight1~19_combout\ : std_logic;
SIGNAL \Selector31~1_combout\ : std_logic;
SIGNAL \Selector31~8_combout\ : std_logic;
SIGNAL \vAluRes~1_RESYN1062_BDD1063\ : std_logic;
SIGNAL \vAluRes~1_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[1]~0_combout\ : std_logic;
SIGNAL \RegFile[15][1]~q\ : std_logic;
SIGNAL \RegFile[14][1]~feeder_combout\ : std_logic;
SIGNAL \RegFile[14][1]~q\ : std_logic;
SIGNAL \RegFile[13][1]~feeder_combout\ : std_logic;
SIGNAL \RegFile[13][1]~q\ : std_logic;
SIGNAL \RegFile[9][1]~q\ : std_logic;
SIGNAL \RegFile[10][1]~q\ : std_logic;
SIGNAL \RegFile[11][1]~q\ : std_logic;
SIGNAL \RegFile[8][1]~feeder_combout\ : std_logic;
SIGNAL \RegFile[8][1]~q\ : std_logic;
SIGNAL \Mux121~14_combout\ : std_logic;
SIGNAL \RegFile[12][1]~feeder_combout\ : std_logic;
SIGNAL \RegFile[12][1]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux121~1_combout\ : std_logic;
SIGNAL \RegFile[23][1]~q\ : std_logic;
SIGNAL \RegFile[21][1]~q\ : std_logic;
SIGNAL \RegFile[22][1]~q\ : std_logic;
SIGNAL \RegFile[19][1]~q\ : std_logic;
SIGNAL \RegFile[17][1]~q\ : std_logic;
SIGNAL \RegFile[18][1]~feeder_combout\ : std_logic;
SIGNAL \RegFile[18][1]~q\ : std_logic;
SIGNAL \RegFile[16][1]~q\ : std_logic;
SIGNAL \Mux121~18_combout\ : std_logic;
SIGNAL \RegFile[20][1]~q\ : std_logic;
SIGNAL \Mux121~5_combout\ : std_logic;
SIGNAL \RegFile[29][1]~q\ : std_logic;
SIGNAL \RegFile[31][1]~feeder_combout\ : std_logic;
SIGNAL \RegFile[31][1]~q\ : std_logic;
SIGNAL \RegFile[30][1]~q\ : std_logic;
SIGNAL \RegFile[27][1]~feeder_combout\ : std_logic;
SIGNAL \RegFile[27][1]~q\ : std_logic;
SIGNAL \RegFile[26][1]~feeder_combout\ : std_logic;
SIGNAL \RegFile[26][1]~q\ : std_logic;
SIGNAL \RegFile[25][1]~q\ : std_logic;
SIGNAL \RegFile[24][1]~feeder_combout\ : std_logic;
SIGNAL \RegFile[24][1]~q\ : std_logic;
SIGNAL \Mux121~22_combout\ : std_logic;
SIGNAL \RegFile[28][1]~feeder_combout\ : std_logic;
SIGNAL \RegFile[28][1]~q\ : std_logic;
SIGNAL \Mux121~9_combout\ : std_logic;
SIGNAL \RegFile[3][1]~q\ : std_logic;
SIGNAL \RegFile[2][1]~q\ : std_logic;
SIGNAL \RegFile[7][1]~q\ : std_logic;
SIGNAL \RegFile[5][1]~feeder_combout\ : std_logic;
SIGNAL \RegFile[5][1]~q\ : std_logic;
SIGNAL \RegFile[4][1]~q\ : std_logic;
SIGNAL \RegFile[6][1]~q\ : std_logic;
SIGNAL \Mux121~0_combout\ : std_logic;
SIGNAL \RegFile[1][1]~feeder_combout\ : std_logic;
SIGNAL \RegFile[1][1]~q\ : std_logic;
SIGNAL \Mux121~26_combout\ : std_logic;
SIGNAL \Mux121~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[1]~17_combout\ : std_logic;
SIGNAL \Selector18~0_combout\ : std_logic;
SIGNAL \Selector18~1_RTM0433_combout\ : std_logic;
SIGNAL \Selector18~1_OTERM431\ : std_logic;
SIGNAL \Selector18~2_combout\ : std_logic;
SIGNAL \ShiftLeft0~21_combout\ : std_logic;
SIGNAL \ShiftRight1~53_combout\ : std_logic;
SIGNAL \Selector18~3_combout\ : std_logic;
SIGNAL \Selector18~4_combout\ : std_logic;
SIGNAL \Add3~57_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[14]~0_combout\ : std_logic;
SIGNAL \Mux76~14_combout\ : std_logic;
SIGNAL \Mux76~1_combout\ : std_logic;
SIGNAL \Mux76~22_combout\ : std_logic;
SIGNAL \Mux76~9_combout\ : std_logic;
SIGNAL \Mux76~18_combout\ : std_logic;
SIGNAL \Mux76~5_combout\ : std_logic;
SIGNAL \Mux76~0_combout\ : std_logic;
SIGNAL \RegFile[1][14]~q\ : std_logic;
SIGNAL \Mux76~26_combout\ : std_logic;
SIGNAL \Mux76~13_combout\ : std_logic;
SIGNAL \Mux240~0_combout\ : std_logic;
SIGNAL \ShiftLeft0~24_combout\ : std_logic;
SIGNAL \ShiftLeft0~24_OTERM293\ : std_logic;
SIGNAL \ShiftLeft0~33_combout\ : std_logic;
SIGNAL \Selector12~0_combout\ : std_logic;
SIGNAL \ShiftRight1~39_combout\ : std_logic;
SIGNAL \Selector12~1_combout\ : std_logic;
SIGNAL \Selector12~5_combout\ : std_logic;
SIGNAL \Add3~81_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[20]~0_combout\ : std_logic;
SIGNAL \Mux70~0_combout\ : std_logic;
SIGNAL \RegFile[1][20]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux70~26_combout\ : std_logic;
SIGNAL \RegFile[14][20]~q\ : std_logic;
SIGNAL \Mux70~14_combout\ : std_logic;
SIGNAL \Mux70~1_combout\ : std_logic;
SIGNAL \Mux70~22_combout\ : std_logic;
SIGNAL \Mux70~9_combout\ : std_logic;
SIGNAL \RegFile[18][20]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux70~18_combout\ : std_logic;
SIGNAL \Mux70~5_combout\ : std_logic;
SIGNAL \Mux70~13_combout\ : std_logic;
SIGNAL \Mux234~0_combout\ : std_logic;
SIGNAL \ShiftLeft0~36_combout\ : std_logic;
SIGNAL \ShiftLeft0~36_OTERM603\ : std_logic;
SIGNAL \ShiftLeft0~45_combout\ : std_logic;
SIGNAL \ShiftLeft0~45_OTERM757\ : std_logic;
SIGNAL \ShiftLeft0~53_combout\ : std_logic;
SIGNAL \ShiftLeft0~53_OTERM765\ : std_logic;
SIGNAL \ShiftLeft0~54_combout\ : std_logic;
SIGNAL \Selector2~0_combout\ : std_logic;
SIGNAL \Selector2~1_combout\ : std_logic;
SIGNAL \Selector2~2_combout\ : std_logic;
SIGNAL \Comb:vJumpAdr[30]~0_RESYN1036_BDD1037\ : std_logic;
SIGNAL \Add3~118\ : std_logic;
SIGNAL \Add3~121_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[30]~0_combout\ : std_logic;
SIGNAL \R.curPC[30]~DUPLICATE_q\ : std_logic;
SIGNAL \Add0~114\ : std_logic;
SIGNAL \Add0~117_sumout\ : std_logic;
SIGNAL \avm_d_readdata[7]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[31]~1_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[31]~2_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[31]~0_combout\ : std_logic;
SIGNAL \RegFile[3][31]~q\ : std_logic;
SIGNAL \RegFile[2][31]~q\ : std_logic;
SIGNAL \RegFile[7][31]~q\ : std_logic;
SIGNAL \RegFile[5][31]~q\ : std_logic;
SIGNAL \RegFile[4][31]~feeder_combout\ : std_logic;
SIGNAL \RegFile[4][31]~q\ : std_logic;
SIGNAL \RegFile[6][31]~q\ : std_logic;
SIGNAL \Mux91~0_combout\ : std_logic;
SIGNAL \RegFile[1][31]~feeder_combout\ : std_logic;
SIGNAL \RegFile[1][31]~q\ : std_logic;
SIGNAL \Mux91~26_combout\ : std_logic;
SIGNAL \RegFile[13][31]~q\ : std_logic;
SIGNAL \RegFile[15][31]~q\ : std_logic;
SIGNAL \RegFile[14][31]~feeder_combout\ : std_logic;
SIGNAL \RegFile[14][31]~q\ : std_logic;
SIGNAL \RegFile[9][31]~q\ : std_logic;
SIGNAL \RegFile[11][31]~q\ : std_logic;
SIGNAL \RegFile[10][31]~feeder_combout\ : std_logic;
SIGNAL \RegFile[10][31]~q\ : std_logic;
SIGNAL \RegFile[8][31]~q\ : std_logic;
SIGNAL \Mux91~14_combout\ : std_logic;
SIGNAL \RegFile[12][31]~feeder_combout\ : std_logic;
SIGNAL \RegFile[12][31]~q\ : std_logic;
SIGNAL \Mux91~1_combout\ : std_logic;
SIGNAL \RegFile[29][31]~q\ : std_logic;
SIGNAL \RegFile[30][31]~q\ : std_logic;
SIGNAL \RegFile[31][31]~q\ : std_logic;
SIGNAL \RegFile[25][31]~q\ : std_logic;
SIGNAL \RegFile[27][31]~q\ : std_logic;
SIGNAL \RegFile[26][31]~q\ : std_logic;
SIGNAL \RegFile[24][31]~feeder_combout\ : std_logic;
SIGNAL \RegFile[24][31]~q\ : std_logic;
SIGNAL \Mux91~22_combout\ : std_logic;
SIGNAL \RegFile[28][31]~feeder_combout\ : std_logic;
SIGNAL \RegFile[28][31]~q\ : std_logic;
SIGNAL \Mux91~9_combout\ : std_logic;
SIGNAL \RegFile[21][31]~q\ : std_logic;
SIGNAL \RegFile[23][31]~q\ : std_logic;
SIGNAL \RegFile[22][31]~feeder_combout\ : std_logic;
SIGNAL \RegFile[22][31]~q\ : std_logic;
SIGNAL \RegFile[17][31]~q\ : std_logic;
SIGNAL \RegFile[18][31]~feeder_combout\ : std_logic;
SIGNAL \RegFile[18][31]~q\ : std_logic;
SIGNAL \RegFile[19][31]~feeder_combout\ : std_logic;
SIGNAL \RegFile[19][31]~q\ : std_logic;
SIGNAL \RegFile[16][31]~feeder_combout\ : std_logic;
SIGNAL \RegFile[16][31]~q\ : std_logic;
SIGNAL \Mux91~18_combout\ : std_logic;
SIGNAL \RegFile[20][31]~feeder_combout\ : std_logic;
SIGNAL \RegFile[20][31]~q\ : std_logic;
SIGNAL \Mux91~5_combout\ : std_logic;
SIGNAL \Mux91~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[31]~29_combout\ : std_logic;
SIGNAL \Add2~125_sumout\ : std_logic;
SIGNAL \Selector1~3_combout\ : std_logic;
SIGNAL \vAluRes~30_combout\ : std_logic;
SIGNAL \vAluRes~29_combout\ : std_logic;
SIGNAL \Add3~122\ : std_logic;
SIGNAL \Add3~125_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[31]~0_combout\ : std_logic;
SIGNAL \R.curPC[31]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux59~0_combout\ : std_logic;
SIGNAL \Mux59~26_combout\ : std_logic;
SIGNAL \RegFile[18][31]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux59~18_combout\ : std_logic;
SIGNAL \Mux59~5_combout\ : std_logic;
SIGNAL \Mux59~14_combout\ : std_logic;
SIGNAL \Mux59~1_combout\ : std_logic;
SIGNAL \Mux59~22_combout\ : std_logic;
SIGNAL \Mux59~9_combout\ : std_logic;
SIGNAL \Mux59~13_combout\ : std_logic;
SIGNAL \Mux223~0_combout\ : std_logic;
SIGNAL \ShiftRight1~48_combout\ : std_logic;
SIGNAL \Selector22~0_OTERM475_OTERM747\ : std_logic;
SIGNAL \ShiftRight0~11_combout\ : std_logic;
SIGNAL \Selector22~0_OTERM475_OTERM749\ : std_logic;
SIGNAL \Selector22~0_RTM0477_combout\ : std_logic;
SIGNAL \ShiftLeft0~46_combout\ : std_logic;
SIGNAL \Selector6~0_combout\ : std_logic;
SIGNAL \ShiftLeft0~44_combout\ : std_logic;
SIGNAL \Selector6~1_combout\ : std_logic;
SIGNAL \Selector6~2_combout\ : std_logic;
SIGNAL \vAluRes~28_combout\ : std_logic;
SIGNAL \Add3~105_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[26]~0_combout\ : std_logic;
SIGNAL \Add0~98\ : std_logic;
SIGNAL \Add0~101_sumout\ : std_logic;
SIGNAL \avm_d_readdata[3]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[27]~1_combout\ : std_logic;
SIGNAL \R.aluRes[27]~DUPLICATE_q\ : std_logic;
SIGNAL \Comb:vRegWriteData[27]~3_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[27]~2_RESYN1108_BDD1109\ : std_logic;
SIGNAL \Comb:vRegWriteData[27]~2_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[27]~0_combout\ : std_logic;
SIGNAL \RegFile[29][27]~q\ : std_logic;
SIGNAL \RegFile[26][27]~q\ : std_logic;
SIGNAL \Mux95~22_combout\ : std_logic;
SIGNAL \Mux95~9_combout\ : std_logic;
SIGNAL \Mux95~0_combout\ : std_logic;
SIGNAL \Mux95~26_combout\ : std_logic;
SIGNAL \Mux95~18_combout\ : std_logic;
SIGNAL \Mux95~5_combout\ : std_logic;
SIGNAL \Mux95~14_combout\ : std_logic;
SIGNAL \Mux95~1_combout\ : std_logic;
SIGNAL \Mux95~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[27]~24_combout\ : std_logic;
SIGNAL \Add1~109_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[27]~0_RESYN1030_BDD1031\ : std_logic;
SIGNAL \Add3~109_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[27]~0_combout\ : std_logic;
SIGNAL \Add0~102\ : std_logic;
SIGNAL \Add0~105_sumout\ : std_logic;
SIGNAL \avm_d_readdata[4]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[28]~1_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[28]~2_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[28]~0_combout\ : std_logic;
SIGNAL \RegFile[13][28]~q\ : std_logic;
SIGNAL \RegFile[15][28]~q\ : std_logic;
SIGNAL \RegFile[14][28]~feeder_combout\ : std_logic;
SIGNAL \RegFile[14][28]~q\ : std_logic;
SIGNAL \RegFile[11][28]~q\ : std_logic;
SIGNAL \RegFile[9][28]~feeder_combout\ : std_logic;
SIGNAL \RegFile[9][28]~q\ : std_logic;
SIGNAL \RegFile[10][28]~feeder_combout\ : std_logic;
SIGNAL \RegFile[10][28]~q\ : std_logic;
SIGNAL \RegFile[8][28]~feeder_combout\ : std_logic;
SIGNAL \RegFile[8][28]~q\ : std_logic;
SIGNAL \Mux94~14_combout\ : std_logic;
SIGNAL \RegFile[12][28]~feeder_combout\ : std_logic;
SIGNAL \RegFile[12][28]~q\ : std_logic;
SIGNAL \Mux94~1_combout\ : std_logic;
SIGNAL \RegFile[31][28]~q\ : std_logic;
SIGNAL \RegFile[29][28]~q\ : std_logic;
SIGNAL \RegFile[30][28]~q\ : std_logic;
SIGNAL \RegFile[27][28]~q\ : std_logic;
SIGNAL \RegFile[25][28]~q\ : std_logic;
SIGNAL \RegFile[26][28]~feeder_combout\ : std_logic;
SIGNAL \RegFile[26][28]~q\ : std_logic;
SIGNAL \RegFile[24][28]~feeder_combout\ : std_logic;
SIGNAL \RegFile[24][28]~q\ : std_logic;
SIGNAL \Mux94~22_combout\ : std_logic;
SIGNAL \RegFile[28][28]~feeder_combout\ : std_logic;
SIGNAL \RegFile[28][28]~q\ : std_logic;
SIGNAL \Mux94~9_combout\ : std_logic;
SIGNAL \RegFile[3][28]~q\ : std_logic;
SIGNAL \RegFile[2][28]~q\ : std_logic;
SIGNAL \RegFile[5][28]~q\ : std_logic;
SIGNAL \RegFile[4][28]~feeder_combout\ : std_logic;
SIGNAL \RegFile[4][28]~q\ : std_logic;
SIGNAL \RegFile[7][28]~q\ : std_logic;
SIGNAL \RegFile[6][28]~q\ : std_logic;
SIGNAL \Mux94~0_combout\ : std_logic;
SIGNAL \RegFile[1][28]~feeder_combout\ : std_logic;
SIGNAL \RegFile[1][28]~q\ : std_logic;
SIGNAL \Mux94~26_combout\ : std_logic;
SIGNAL \RegFile[23][28]~q\ : std_logic;
SIGNAL \RegFile[21][28]~feeder_combout\ : std_logic;
SIGNAL \RegFile[21][28]~q\ : std_logic;
SIGNAL \RegFile[22][28]~q\ : std_logic;
SIGNAL \RegFile[19][28]~q\ : std_logic;
SIGNAL \RegFile[17][28]~feeder_combout\ : std_logic;
SIGNAL \RegFile[17][28]~q\ : std_logic;
SIGNAL \RegFile[18][28]~feeder_combout\ : std_logic;
SIGNAL \RegFile[18][28]~q\ : std_logic;
SIGNAL \RegFile[16][28]~feeder_combout\ : std_logic;
SIGNAL \RegFile[16][28]~q\ : std_logic;
SIGNAL \Mux94~18_combout\ : std_logic;
SIGNAL \RegFile[20][28]~q\ : std_logic;
SIGNAL \Mux94~5_combout\ : std_logic;
SIGNAL \Mux94~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[28]~23_combout\ : std_logic;
SIGNAL \Add1~113_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[28]~0_RESYN1032_BDD1033\ : std_logic;
SIGNAL \Add3~113_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[28]~0_combout\ : std_logic;
SIGNAL \Mux62~14_combout\ : std_logic;
SIGNAL \Mux62~1_combout\ : std_logic;
SIGNAL \RegFile[6][28]~DUPLICATE_q\ : std_logic;
SIGNAL \Mux62~0_combout\ : std_logic;
SIGNAL \Mux62~26_combout\ : std_logic;
SIGNAL \Mux62~22_combout\ : std_logic;
SIGNAL \Mux62~9_combout\ : std_logic;
SIGNAL \Mux62~18_combout\ : std_logic;
SIGNAL \Mux62~5_combout\ : std_logic;
SIGNAL \Mux62~13_combout\ : std_logic;
SIGNAL \Mux226~0_combout\ : std_logic;
SIGNAL \ShiftRight1~27_combout\ : std_logic;
SIGNAL \ShiftRight1~27_OTERM19\ : std_logic;
SIGNAL \ShiftRight1~29_combout\ : std_logic;
SIGNAL \Add1~9_sumout\ : std_logic;
SIGNAL \Selector30~0_combout\ : std_logic;
SIGNAL \ShiftRight1~20_combout\ : std_logic;
SIGNAL \ShiftRight1~24_combout\ : std_logic;
SIGNAL \Selector30~1_RTM0405_combout\ : std_logic;
SIGNAL \Selector30~1_OTERM403\ : std_logic;
SIGNAL \Selector30~2_combout\ : std_logic;
SIGNAL \Add2~9_sumout\ : std_logic;
SIGNAL \Selector30~3_combout\ : std_logic;
SIGNAL \Selector30~4_combout\ : std_logic;
SIGNAL \vAluRes~2_RESYN1064_BDD1065\ : std_logic;
SIGNAL \vAluRes~2_combout\ : std_logic;
SIGNAL \Add3~9_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[2]~0_combout\ : std_logic;
SIGNAL \Add0~1_sumout\ : std_logic;
SIGNAL \R.regWriteData[2]~feeder_combout\ : std_logic;
SIGNAL \avm_d_readdata[26]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[2]~0_RESYN1082_BDD1083\ : std_logic;
SIGNAL \Comb:vRegWriteData[2]~0_combout\ : std_logic;
SIGNAL \RegFile[2][2]~q\ : std_logic;
SIGNAL \Mux120~0_combout\ : std_logic;
SIGNAL \Mux120~26_combout\ : std_logic;
SIGNAL \RegFile[14][2]~q\ : std_logic;
SIGNAL \Mux120~14_combout\ : std_logic;
SIGNAL \Mux120~1_combout\ : std_logic;
SIGNAL \Mux120~18_combout\ : std_logic;
SIGNAL \Mux120~5_combout\ : std_logic;
SIGNAL \Mux120~22_combout\ : std_logic;
SIGNAL \Mux120~9_combout\ : std_logic;
SIGNAL \Mux120~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[2]~19_combout\ : std_logic;
SIGNAL \Selector32~3_combout\ : std_logic;
SIGNAL \Selector32~3_OTERM379\ : std_logic;
SIGNAL \Selector31~2_RTM0401_combout\ : std_logic;
SIGNAL \Selector31~2_OTERM399\ : std_logic;
SIGNAL \Selector31~3_combout\ : std_logic;
SIGNAL \Selector31~4_combout\ : std_logic;
SIGNAL \Add3~5_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[1]~0_combout\ : std_logic;
SIGNAL \Mux89~0_combout\ : std_logic;
SIGNAL \Mux89~26_combout\ : std_logic;
SIGNAL \Mux89~22_combout\ : std_logic;
SIGNAL \Mux89~9_combout\ : std_logic;
SIGNAL \Mux89~14_combout\ : std_logic;
SIGNAL \RegFile[12][1]~q\ : std_logic;
SIGNAL \Mux89~1_combout\ : std_logic;
SIGNAL \Mux89~18_combout\ : std_logic;
SIGNAL \Mux89~5_combout\ : std_logic;
SIGNAL \Mux89~13_combout\ : std_logic;
SIGNAL \Mux253~0_combout\ : std_logic;
SIGNAL \ShiftLeft0~5_combout\ : std_logic;
SIGNAL \ShiftLeft0~5_OTERM203\ : std_logic;
SIGNAL \Selector28~1_RTM0389_combout\ : std_logic;
SIGNAL \Selector28~1_OTERM387\ : std_logic;
SIGNAL \Selector28~2_combout\ : std_logic;
SIGNAL \ShiftRight1~6_combout\ : std_logic;
SIGNAL \ShiftRight1~6_OTERM197\ : std_logic;
SIGNAL \ShiftRight1~40_combout\ : std_logic;
SIGNAL \ShiftRight0~6_combout\ : std_logic;
SIGNAL \Selector28~3_combout\ : std_logic;
SIGNAL \Add2~17_sumout\ : std_logic;
SIGNAL \Add1~17_sumout\ : std_logic;
SIGNAL \Selector28~0_combout\ : std_logic;
SIGNAL \Selector28~4_combout\ : std_logic;
SIGNAL \R.aluRes[4]~DUPLICATE_q\ : std_logic;
SIGNAL \vAluRes~4_RESYN1068_BDD1069\ : std_logic;
SIGNAL \vAluRes~4_combout\ : std_logic;
SIGNAL \Add3~17_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[4]~0_combout\ : std_logic;
SIGNAL \Add0~9_sumout\ : std_logic;
SIGNAL \R.regWriteData[4]~feeder_combout\ : std_logic;
SIGNAL \avm_d_readdata[28]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[4]~0_RESYN1090_BDD1091\ : std_logic;
SIGNAL \Comb:vRegWriteData[4]~0_combout\ : std_logic;
SIGNAL \RegFile[23][4]~feeder_combout\ : std_logic;
SIGNAL \RegFile[23][4]~q\ : std_logic;
SIGNAL \Mux118~18_combout\ : std_logic;
SIGNAL \Mux118~5_combout\ : std_logic;
SIGNAL \Mux118~14_combout\ : std_logic;
SIGNAL \Mux118~1_combout\ : std_logic;
SIGNAL \Mux118~0_combout\ : std_logic;
SIGNAL \Mux118~26_combout\ : std_logic;
SIGNAL \Mux118~22_combout\ : std_logic;
SIGNAL \Mux118~9_combout\ : std_logic;
SIGNAL \Mux118~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[4]~20_combout\ : std_logic;
SIGNAL \Selector12~2_combout\ : std_logic;
SIGNAL \Selector12~2_OTERM395\ : std_logic;
SIGNAL \Selector11~2_combout\ : std_logic;
SIGNAL \Selector11~3_combout\ : std_logic;
SIGNAL \Selector11~4_combout\ : std_logic;
SIGNAL \Selector11~5_combout\ : std_logic;
SIGNAL \Add3~85_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[21]~0_combout\ : std_logic;
SIGNAL \R.curPC[21]~DUPLICATE_q\ : std_logic;
SIGNAL \Add0~77_sumout\ : std_logic;
SIGNAL \R.regWriteData[21]~feeder_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[21]~1_RESYN1130_BDD1131\ : std_logic;
SIGNAL \avm_d_readdata[13]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[21]~1_RESYN1126_BDD1127\ : std_logic;
SIGNAL \Comb:vRegWriteData[21]~1_RESYN1128_BDD1129\ : std_logic;
SIGNAL \Comb:vRegWriteData[21]~1_combout\ : std_logic;
SIGNAL \RegFile[3][21]~q\ : std_logic;
SIGNAL \Mux101~0_combout\ : std_logic;
SIGNAL \Mux101~26_combout\ : std_logic;
SIGNAL \Mux101~14_combout\ : std_logic;
SIGNAL \Mux101~1_combout\ : std_logic;
SIGNAL \Mux101~18_combout\ : std_logic;
SIGNAL \Mux101~5_combout\ : std_logic;
SIGNAL \Mux101~22_combout\ : std_logic;
SIGNAL \Mux101~9_combout\ : std_logic;
SIGNAL \Mux101~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[21]~0_combout\ : std_logic;
SIGNAL \Add1~86\ : std_logic;
SIGNAL \Add1~89_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[22]~0_RESYN1028_BDD1029\ : std_logic;
SIGNAL \Add3~89_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[22]~0_combout\ : std_logic;
SIGNAL \Add0~81_sumout\ : std_logic;
SIGNAL \Comb:vRegWriteData[22]~3_combout\ : std_logic;
SIGNAL \avm_d_readdata[14]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[22]~2_RESYN1112_BDD1113\ : std_logic;
SIGNAL \Comb:vRegWriteData[22]~2_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[22]~1_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[22]~0_combout\ : std_logic;
SIGNAL \RegFile[31][22]~q\ : std_logic;
SIGNAL \Mux100~22_combout\ : std_logic;
SIGNAL \Mux100~9_combout\ : std_logic;
SIGNAL \Mux100~14_combout\ : std_logic;
SIGNAL \Mux100~1_combout\ : std_logic;
SIGNAL \Mux100~18_combout\ : std_logic;
SIGNAL \Mux100~5_combout\ : std_logic;
SIGNAL \Mux100~0_combout\ : std_logic;
SIGNAL \Mux100~26_combout\ : std_logic;
SIGNAL \Mux100~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[22]~28_combout\ : std_logic;
SIGNAL \Add1~90\ : std_logic;
SIGNAL \Add1~93_sumout\ : std_logic;
SIGNAL \ShiftRight0~12_combout\ : std_logic;
SIGNAL \ShiftLeft0~39_combout\ : std_logic;
SIGNAL \Selector9~0_combout\ : std_logic;
SIGNAL \Selector9~1_combout\ : std_logic;
SIGNAL \Add2~93_sumout\ : std_logic;
SIGNAL \Selector9~3_combout\ : std_logic;
SIGNAL \LessThan1~30_combout\ : std_logic;
SIGNAL \LessThan1~30_OTERM43\ : std_logic;
SIGNAL \Selector9~2_combout\ : std_logic;
SIGNAL \Selector9~4_combout\ : std_logic;
SIGNAL \Selector9~5_combout\ : std_logic;
SIGNAL \Add3~93_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[23]~0_combout\ : std_logic;
SIGNAL \Add0~85_sumout\ : std_logic;
SIGNAL \avm_d_readdata[15]~input_o\ : std_logic;
SIGNAL \Comb:vRegWriteData[23]~1_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[23]~3_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[23]~2_RESYN1114_BDD1115\ : std_logic;
SIGNAL \Comb:vRegWriteData[23]~2_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[23]~0_combout\ : std_logic;
SIGNAL \RegFile[15][23]~q\ : std_logic;
SIGNAL \Mux99~14_combout\ : std_logic;
SIGNAL \Mux99~1_combout\ : std_logic;
SIGNAL \RegFile[16][23]~q\ : std_logic;
SIGNAL \Mux99~18_combout\ : std_logic;
SIGNAL \Mux99~5_combout\ : std_logic;
SIGNAL \Mux99~22_combout\ : std_logic;
SIGNAL \Mux99~9_combout\ : std_logic;
SIGNAL \Mux99~0_combout\ : std_logic;
SIGNAL \Mux99~26_combout\ : std_logic;
SIGNAL \Mux99~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[23]~27_combout\ : std_logic;
SIGNAL \LessThan1~29_combout\ : std_logic;
SIGNAL \LessThan1~29_OTERM47\ : std_logic;
SIGNAL \LessThan1~28_RTM053_combout\ : std_logic;
SIGNAL \LessThan1~28_OTERM51\ : std_logic;
SIGNAL \LessThan1~33_combout\ : std_logic;
SIGNAL \LessThan1~34_combout\ : std_logic;
SIGNAL \LessThan1~34_OTERM55\ : std_logic;
SIGNAL \LessThan1~35_combout\ : std_logic;
SIGNAL \LessThan1~36_combout\ : std_logic;
SIGNAL \LessThan1~38_combout\ : std_logic;
SIGNAL \LessThan1~37_combout\ : std_logic;
SIGNAL \Mux20~0_combout\ : std_logic;
SIGNAL \Mux20~1_combout\ : std_logic;
SIGNAL \R.aluOp.ALUOpSLTU_OTERM571\ : std_logic;
SIGNAL \R.aluOp.ALUOpSLTU~q\ : std_logic;
SIGNAL \Mux221~0_combout\ : std_logic;
SIGNAL \Mux19~0_combout\ : std_logic;
SIGNAL \R.aluOp.ALUOpSLT_OTERM573\ : std_logic;
SIGNAL \R.aluOp.ALUOpSLT~q\ : std_logic;
SIGNAL \Selector32~0_combout\ : std_logic;
SIGNAL \LessThan1~32_combout\ : std_logic;
SIGNAL \LessThan1~0_RTM0345_combout\ : std_logic;
SIGNAL \LessThan1~0_OTERM343\ : std_logic;
SIGNAL \LessThan1~2_RTM0333_combout\ : std_logic;
SIGNAL \LessThan1~2_OTERM331\ : std_logic;
SIGNAL \LessThan1~1_RTM0339_combout\ : std_logic;
SIGNAL \LessThan1~1_OTERM337\ : std_logic;
SIGNAL \LessThan1~3_RTM0327_combout\ : std_logic;
SIGNAL \LessThan1~3_OTERM325\ : std_logic;
SIGNAL \LessThan1~25_combout\ : std_logic;
SIGNAL \LessThan1~25_OTERM317\ : std_logic;
SIGNAL \LessThan1~24_combout\ : std_logic;
SIGNAL \LessThan1~24_OTERM329\ : std_logic;
SIGNAL \LessThan1~26_combout\ : std_logic;
SIGNAL \LessThan1~4_combout\ : std_logic;
SIGNAL \LessThan1~4_OTERM319\ : std_logic;
SIGNAL \LessThan1~5_RTM0315_combout\ : std_logic;
SIGNAL \LessThan1~5_OTERM313\ : std_logic;
SIGNAL \LessThan1~6_combout\ : std_logic;
SIGNAL \LessThan1~20_combout\ : std_logic;
SIGNAL \LessThan1~20_OTERM341\ : std_logic;
SIGNAL \LessThan1~22_combout\ : std_logic;
SIGNAL \LessThan1~22_OTERM347\ : std_logic;
SIGNAL \LessThan1~21_combout\ : std_logic;
SIGNAL \LessThan1~21_OTERM335\ : std_logic;
SIGNAL \LessThan1~23_combout\ : std_logic;
SIGNAL \LessThan1~18_RTM0323_combout\ : std_logic;
SIGNAL \LessThan1~18_OTERM321\ : std_logic;
SIGNAL \LessThan1~19_combout\ : std_logic;
SIGNAL \LessThan1~7_RTM0309_combout\ : std_logic;
SIGNAL \LessThan1~7_OTERM307\ : std_logic;
SIGNAL \LessThan1~10_RTM0215_combout\ : std_logic;
SIGNAL \LessThan1~10_OTERM213\ : std_logic;
SIGNAL \LessThan1~8_RTM0303_combout\ : std_logic;
SIGNAL \LessThan1~8_OTERM301\ : std_logic;
SIGNAL \LessThan1~9_combout\ : std_logic;
SIGNAL \LessThan1~9_OTERM253\ : std_logic;
SIGNAL \LessThan1~11_combout\ : std_logic;
SIGNAL \LessThan1~11_OTERM217\ : std_logic;
SIGNAL \LessThan1~12_RTM0193_combout\ : std_logic;
SIGNAL \LessThan1~12_OTERM191\ : std_logic;
SIGNAL \LessThan1~13_combout\ : std_logic;
SIGNAL \LessThan1~14_combout\ : std_logic;
SIGNAL \LessThan1~14_OTERM305\ : std_logic;
SIGNAL \LessThan1~15_combout\ : std_logic;
SIGNAL \LessThan1~15_OTERM195\ : std_logic;
SIGNAL \LessThan1~16_combout\ : std_logic;
SIGNAL \LessThan1~16_OTERM311\ : std_logic;
SIGNAL \LessThan1~17_combout\ : std_logic;
SIGNAL \LessThan1~27_combout\ : std_logic;
SIGNAL \Selector32~1_combout\ : std_logic;
SIGNAL \Selector32~8_combout\ : std_logic;
SIGNAL \Comb:vRegWriteData[0]~1_combout\ : std_logic;
SIGNAL \RegFile[3][0]~q\ : std_logic;
SIGNAL \Mux122~0_combout\ : std_logic;
SIGNAL \Mux122~26_combout\ : std_logic;
SIGNAL \Mux122~22_combout\ : std_logic;
SIGNAL \RegFile[28][0]~q\ : std_logic;
SIGNAL \Mux122~9_combout\ : std_logic;
SIGNAL \RegFile[18][0]~q\ : std_logic;
SIGNAL \Mux122~18_combout\ : std_logic;
SIGNAL \Mux122~5_combout\ : std_logic;
SIGNAL \Mux122~14_combout\ : std_logic;
SIGNAL \RegFile[12][0]~q\ : std_logic;
SIGNAL \Mux122~1_combout\ : std_logic;
SIGNAL \Mux122~13_combout\ : std_logic;
SIGNAL \NxR.aluData2[0]~16_combout\ : std_logic;
SIGNAL \Add2~1_sumout\ : std_logic;
SIGNAL \Selector32~4_combout\ : std_logic;
SIGNAL \Selector32~4_OTERM397\ : std_logic;
SIGNAL \Selector32~7_RESYN1056_BDD1057\ : std_logic;
SIGNAL \Selector32~7_RESYN1058_BDD1059\ : std_logic;
SIGNAL \ShiftRight1~5_combout\ : std_logic;
SIGNAL \ShiftRight1~5_OTERM219\ : std_logic;
SIGNAL \ShiftRight1~9_combout\ : std_logic;
SIGNAL \Selector32~7_RESYN1060_BDD1061\ : std_logic;
SIGNAL \Selector32~2_combout\ : std_logic;
SIGNAL \Selector32~7_combout\ : std_logic;
SIGNAL \Add3~1_sumout\ : std_logic;
SIGNAL \Comb:vJumpAdr[0]~0_combout\ : std_logic;
SIGNAL \R.curPC[0]~DUPLICATE_q\ : std_logic;
SIGNAL \R.curPC[29]~DUPLICATE_q\ : std_logic;
SIGNAL \vAluRes~9_combout\ : std_logic;
SIGNAL \vAluRes~11_combout\ : std_logic;
SIGNAL \vAluRes~12_combout\ : std_logic;
SIGNAL \Selector16~4_combout\ : std_logic;
SIGNAL \vAluRes~13_combout\ : std_logic;
SIGNAL \Selector15~1_combout\ : std_logic;
SIGNAL \vAluRes~14_combout\ : std_logic;
SIGNAL \vAluRes~15_combout\ : std_logic;
SIGNAL \vAluRes~16_combout\ : std_logic;
SIGNAL \vAluRes~18_combout\ : std_logic;
SIGNAL \vAluRes~20_combout\ : std_logic;
SIGNAL \vAluRes~21_combout\ : std_logic;
SIGNAL \vAluRes~22_combout\ : std_logic;
SIGNAL \vAluRes~23_combout\ : std_logic;
SIGNAL \Mux221~1_combout\ : std_logic;
SIGNAL \NxR~6_combout\ : std_logic;
SIGNAL \R.memWrite~q\ : std_logic;
SIGNAL \Mux194~0_combout\ : std_logic;
SIGNAL \Mux193~0_combout\ : std_logic;
SIGNAL \Mux192~0_combout\ : std_logic;
SIGNAL \Mux191~0_combout\ : std_logic;
SIGNAL \Mux190~0_combout\ : std_logic;
SIGNAL \Mux189~0_combout\ : std_logic;
SIGNAL \Mux188~0_combout\ : std_logic;
SIGNAL \Mux187~0_combout\ : std_logic;
SIGNAL \Mux202~0_combout\ : std_logic;
SIGNAL \Mux201~0_combout\ : std_logic;
SIGNAL \Mux200~0_combout\ : std_logic;
SIGNAL \Mux199~0_combout\ : std_logic;
SIGNAL \Mux198~0_combout\ : std_logic;
SIGNAL \Mux197~0_combout\ : std_logic;
SIGNAL \Mux196~0_combout\ : std_logic;
SIGNAL \Mux195~0_combout\ : std_logic;
SIGNAL \Mux210~0_combout\ : std_logic;
SIGNAL \Mux209~0_combout\ : std_logic;
SIGNAL \Mux208~0_combout\ : std_logic;
SIGNAL \Mux207~0_combout\ : std_logic;
SIGNAL \Mux206~0_combout\ : std_logic;
SIGNAL \Mux205~0_combout\ : std_logic;
SIGNAL \Mux204~0_combout\ : std_logic;
SIGNAL \Mux203~0_combout\ : std_logic;
SIGNAL \Mux218~0_combout\ : std_logic;
SIGNAL \Mux217~0_combout\ : std_logic;
SIGNAL \Mux216~0_combout\ : std_logic;
SIGNAL \Mux215~0_combout\ : std_logic;
SIGNAL \Mux214~0_combout\ : std_logic;
SIGNAL \Mux213~0_combout\ : std_logic;
SIGNAL \Mux212~0_combout\ : std_logic;
SIGNAL \Mux211~0_combout\ : std_logic;
SIGNAL \NxR~7_combout\ : std_logic;
SIGNAL \R.memRead~q\ : std_logic;
SIGNAL \R.curPC\ : std_logic_vector(31 DOWNTO 0);
SIGNAL \R.regWriteData\ : std_logic_vector(31 DOWNTO 0);
SIGNAL \R.aluData1\ : std_logic_vector(31 DOWNTO 0);
SIGNAL \R.aluData2\ : std_logic_vector(31 DOWNTO 0);
SIGNAL \R.aluRes\ : std_logic_vector(31 DOWNTO 0);
SIGNAL \R.curInst\ : std_logic_vector(31 DOWNTO 0);
SIGNAL \R.statusReg\ : std_logic_vector(31 DOWNTO 0);
SIGNAL \ALT_INV_Add3~5_sumout\ : std_logic;
SIGNAL \ALT_INV_R.jumpToAdr~q\ : std_logic;
SIGNAL \ALT_INV_Add3~1_sumout\ : std_logic;
SIGNAL \ALT_INV_Mux99~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux99~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux99~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux100~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux100~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux100~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux101~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux101~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux101~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux102~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux102~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux102~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux103~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux103~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux103~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux104~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux104~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux104~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux105~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux105~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux105~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux106~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux106~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux106~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux115~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux115~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux115~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux107~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux107~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux107~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux91~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux91~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux91~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux116~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux116~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux116~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux108~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux108~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux108~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux92~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux92~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux92~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux117~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux117~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux117~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux109~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux109~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux109~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux93~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux93~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux93~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux118~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux118~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux118~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux110~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux110~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux110~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux94~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux94~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux94~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux119~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux119~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux119~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux111~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux111~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux111~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux95~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux95~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux95~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux120~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux120~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux120~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux112~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux112~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux112~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux96~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux96~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux96~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux121~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux121~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux121~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux113~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux113~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux113~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux97~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux97~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux97~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux122~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux122~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux122~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux114~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux114~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux114~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux98~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux98~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux98~1_combout\ : std_logic;
SIGNAL \ALT_INV_Add1~125_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~125_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~121_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~121_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~117_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~117_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~113_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~113_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~109_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~109_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~105_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~105_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~101_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~101_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~97_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~97_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~93_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~93_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~89_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~89_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~85_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~85_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~81_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~81_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~77_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~77_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~73_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~73_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~69_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~69_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~65_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~65_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~61_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~61_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~57_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~57_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~53_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~53_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~49_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~49_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~45_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~45_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~41_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~41_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~37_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~37_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~33_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~33_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~29_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~29_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~25_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~25_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~21_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~21_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~17_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~17_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~13_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~13_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~9_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~9_sumout\ : std_logic;
SIGNAL \ALT_INV_Add1~5_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~5_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~1_sumout\ : std_logic;
SIGNAL \ALT_INV_R.aluCalc~q\ : std_logic;
SIGNAL \ALT_INV_R.curPC\ : std_logic_vector(31 DOWNTO 1);
SIGNAL \ALT_INV_Mux240~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux76~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux76~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR.aluData2[15]~6_combout\ : std_logic;
SIGNAL \ALT_INV_Mux139~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux239~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux75~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux75~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR.aluData2[16]~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux138~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux238~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux74~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux74~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR.aluData2[17]~4_combout\ : std_logic;
SIGNAL \ALT_INV_Mux137~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux237~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux73~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux73~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR.aluData2[18]~3_combout\ : std_logic;
SIGNAL \ALT_INV_Mux136~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux236~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux72~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux72~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR.aluData2[19]~2_combout\ : std_logic;
SIGNAL \ALT_INV_Mux135~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux123~2_combout\ : std_logic;
SIGNAL \ALT_INV_Mux149~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux235~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux71~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux71~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR.aluData2[20]~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux134~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux234~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux70~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux70~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR.aluData2[21]~0_combout\ : std_logic;
SIGNAL \ALT_INV_vAluSrc2~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux133~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux123~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux124~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux233~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux69~13_combout\ : std_logic;
SIGNAL \ALT_INV_R.curInst\ : std_logic_vector(31 DOWNTO 0);
SIGNAL \ALT_INV_Mux69~0_combout\ : std_logic;
SIGNAL \ALT_INV_vAluSrc1~2_combout\ : std_logic;
SIGNAL \ALT_INV_vAluSrc1~1_combout\ : std_logic;
SIGNAL \ALT_INV_vAluSrc2~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux20~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux20~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux26~0_combout\ : std_logic;
SIGNAL \ALT_INV_R.ctrlState.Fetch~q\ : std_logic;
SIGNAL \ALT_INV_Mux12~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR~4_combout\ : std_logic;
SIGNAL \ALT_INV_Mux154~0_combout\ : std_logic;
SIGNAL \ALT_INV_R.ctrlState.ReadReg~q\ : std_logic;
SIGNAL \ALT_INV_NxR~2_combout\ : std_logic;
SIGNAL \ALT_INV_vAluSrc1~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux123~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux53~2_combout\ : std_logic;
SIGNAL \ALT_INV_R.ctrlState.DataAccess1~q\ : std_logic;
SIGNAL \ALT_INV_NxR~0_combout\ : std_logic;
SIGNAL \ALT_INV_Equal2~2_combout\ : std_logic;
SIGNAL \ALT_INV_Equal2~1_combout\ : std_logic;
SIGNAL \ALT_INV_Equal2~0_combout\ : std_logic;
SIGNAL \ALT_INV_R.ctrlState.Trap~q\ : std_logic;
SIGNAL \ALT_INV_R.ctrlState.Wait0~q\ : std_logic;
SIGNAL \ALT_INV_Mux53~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux53~0_combout\ : std_logic;
SIGNAL \ALT_INV_R.ctrlState.DataAccess0~q\ : std_logic;
SIGNAL \ALT_INV_R.ctrlState.Calc~q\ : std_logic;
SIGNAL \ALT_INV_Mux18~0_combout\ : std_logic;
SIGNAL \ALT_INV_vAluRes~30_combout\ : std_logic;
SIGNAL \ALT_INV_vAluRes~29_combout\ : std_logic;
SIGNAL \ALT_INV_vAluRes~28_combout\ : std_logic;
SIGNAL \ALT_INV_vAluRes~27_combout\ : std_logic;
SIGNAL \ALT_INV_vAluRes~26_combout\ : std_logic;
SIGNAL \ALT_INV_vAluRes~25_combout\ : std_logic;
SIGNAL \ALT_INV_Selector7~4_combout\ : std_logic;
SIGNAL \ALT_INV_Selector13~2_combout\ : std_logic;
SIGNAL \ALT_INV_Selector14~4_combout\ : std_logic;
SIGNAL \ALT_INV_Selector15~5_combout\ : std_logic;
SIGNAL \ALT_INV_Selector16~5_combout\ : std_logic;
SIGNAL \ALT_INV_Equal4~2_combout\ : std_logic;
SIGNAL \ALT_INV_Equal4~1_combout\ : std_logic;
SIGNAL \ALT_INV_Equal4~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux99~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][23]~q\ : std_logic;
SIGNAL \ALT_INV_Mux99~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][23]~q\ : std_logic;
SIGNAL \ALT_INV_Mux100~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][22]~q\ : std_logic;
SIGNAL \ALT_INV_Mux100~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][22]~q\ : std_logic;
SIGNAL \ALT_INV_Mux101~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][21]~q\ : std_logic;
SIGNAL \ALT_INV_Mux101~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][21]~q\ : std_logic;
SIGNAL \ALT_INV_Mux102~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][20]~q\ : std_logic;
SIGNAL \ALT_INV_Mux102~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][20]~q\ : std_logic;
SIGNAL \ALT_INV_Mux103~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][19]~q\ : std_logic;
SIGNAL \ALT_INV_Mux103~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][19]~q\ : std_logic;
SIGNAL \ALT_INV_Mux104~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][18]~q\ : std_logic;
SIGNAL \ALT_INV_Mux104~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][18]~q\ : std_logic;
SIGNAL \ALT_INV_Mux105~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][17]~q\ : std_logic;
SIGNAL \ALT_INV_Mux105~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][17]~q\ : std_logic;
SIGNAL \ALT_INV_Mux106~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][16]~q\ : std_logic;
SIGNAL \ALT_INV_Mux106~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][16]~q\ : std_logic;
SIGNAL \ALT_INV_Mux115~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][7]~q\ : std_logic;
SIGNAL \ALT_INV_Mux115~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][7]~q\ : std_logic;
SIGNAL \ALT_INV_Mux107~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][15]~q\ : std_logic;
SIGNAL \ALT_INV_Mux107~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][15]~q\ : std_logic;
SIGNAL \ALT_INV_Mux91~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][31]~q\ : std_logic;
SIGNAL \ALT_INV_Mux91~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][31]~q\ : std_logic;
SIGNAL \ALT_INV_Mux116~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][6]~q\ : std_logic;
SIGNAL \ALT_INV_Mux116~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][6]~q\ : std_logic;
SIGNAL \ALT_INV_Mux108~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][14]~q\ : std_logic;
SIGNAL \ALT_INV_Mux108~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][14]~q\ : std_logic;
SIGNAL \ALT_INV_Mux92~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][30]~q\ : std_logic;
SIGNAL \ALT_INV_Mux92~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][30]~q\ : std_logic;
SIGNAL \ALT_INV_Mux117~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][5]~q\ : std_logic;
SIGNAL \ALT_INV_Mux117~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][5]~q\ : std_logic;
SIGNAL \ALT_INV_Mux109~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][13]~q\ : std_logic;
SIGNAL \ALT_INV_Mux109~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][13]~q\ : std_logic;
SIGNAL \ALT_INV_Mux93~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][29]~q\ : std_logic;
SIGNAL \ALT_INV_Mux93~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][29]~q\ : std_logic;
SIGNAL \ALT_INV_Mux118~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][4]~q\ : std_logic;
SIGNAL \ALT_INV_Mux118~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][4]~q\ : std_logic;
SIGNAL \ALT_INV_Mux110~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][12]~q\ : std_logic;
SIGNAL \ALT_INV_Mux110~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][12]~q\ : std_logic;
SIGNAL \ALT_INV_Mux94~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][28]~q\ : std_logic;
SIGNAL \ALT_INV_Mux94~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][28]~q\ : std_logic;
SIGNAL \ALT_INV_Mux119~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][3]~q\ : std_logic;
SIGNAL \ALT_INV_Mux119~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][3]~q\ : std_logic;
SIGNAL \ALT_INV_Mux111~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][11]~q\ : std_logic;
SIGNAL \ALT_INV_Mux111~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][11]~q\ : std_logic;
SIGNAL \ALT_INV_Mux95~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][27]~q\ : std_logic;
SIGNAL \ALT_INV_Mux95~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][27]~q\ : std_logic;
SIGNAL \ALT_INV_Mux120~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][2]~q\ : std_logic;
SIGNAL \ALT_INV_Mux120~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][2]~q\ : std_logic;
SIGNAL \ALT_INV_Mux112~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][10]~q\ : std_logic;
SIGNAL \ALT_INV_Mux112~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][10]~q\ : std_logic;
SIGNAL \ALT_INV_Mux96~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][26]~q\ : std_logic;
SIGNAL \ALT_INV_Mux96~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][26]~q\ : std_logic;
SIGNAL \ALT_INV_Mux121~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][1]~q\ : std_logic;
SIGNAL \ALT_INV_Mux121~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][1]~q\ : std_logic;
SIGNAL \ALT_INV_Mux113~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][9]~q\ : std_logic;
SIGNAL \ALT_INV_Mux113~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][9]~q\ : std_logic;
SIGNAL \ALT_INV_Mux97~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][25]~q\ : std_logic;
SIGNAL \ALT_INV_Mux97~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][25]~q\ : std_logic;
SIGNAL \ALT_INV_Mux122~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][0]~q\ : std_logic;
SIGNAL \ALT_INV_Mux122~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][0]~q\ : std_logic;
SIGNAL \ALT_INV_Mux114~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][8]~q\ : std_logic;
SIGNAL \ALT_INV_Mux114~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][8]~q\ : std_logic;
SIGNAL \ALT_INV_Mux98~13_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[3][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][24]~q\ : std_logic;
SIGNAL \ALT_INV_Mux98~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][24]~q\ : std_logic;
SIGNAL \ALT_INV_Mux162~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux221~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux222~0_combout\ : std_logic;
SIGNAL \ALT_INV_R.aluRes\ : std_logic_vector(31 DOWNTO 0);
SIGNAL \ALT_INV_Selector1~2_combout\ : std_logic;
SIGNAL \ALT_INV_Selector1~1_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~56_combout\ : std_logic;
SIGNAL \ALT_INV_Selector2~2_combout\ : std_logic;
SIGNAL \ALT_INV_Selector2~1_combout\ : std_logic;
SIGNAL \ALT_INV_Selector2~0_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~54_combout\ : std_logic;
SIGNAL \ALT_INV_Selector3~2_combout\ : std_logic;
SIGNAL \ALT_INV_Selector3~1_combout\ : std_logic;
SIGNAL \ALT_INV_Selector3~0_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~52_combout\ : std_logic;
SIGNAL \ALT_INV_Selector4~1_combout\ : std_logic;
SIGNAL \ALT_INV_Selector4~0_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~50_combout\ : std_logic;
SIGNAL \ALT_INV_Selector20~5_combout\ : std_logic;
SIGNAL \ALT_INV_Selector5~4_combout\ : std_logic;
SIGNAL \ALT_INV_Selector5~3_combout\ : std_logic;
SIGNAL \ALT_INV_Selector5~2_combout\ : std_logic;
SIGNAL \ALT_INV_Selector5~1_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~48_combout\ : std_logic;
SIGNAL \ALT_INV_Selector5~0_combout\ : std_logic;
SIGNAL \ALT_INV_Selector6~2_combout\ : std_logic;
SIGNAL \ALT_INV_Selector6~1_combout\ : std_logic;
SIGNAL \ALT_INV_Selector6~0_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~46_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~44_combout\ : std_logic;
SIGNAL \ALT_INV_Selector7~3_combout\ : std_logic;
SIGNAL \ALT_INV_Selector7~2_combout\ : std_logic;
SIGNAL \ALT_INV_Selector7~1_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~43_combout\ : std_logic;
SIGNAL \ALT_INV_Selector7~0_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~55_combout\ : std_logic;
SIGNAL \ALT_INV_Selector8~4_combout\ : std_logic;
SIGNAL \ALT_INV_Selector8~3_combout\ : std_logic;
SIGNAL \ALT_INV_Selector8~2_combout\ : std_logic;
SIGNAL \ALT_INV_Selector8~1_combout\ : std_logic;
SIGNAL \ALT_INV_Selector8~0_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~41_combout\ : std_logic;
SIGNAL \ALT_INV_Selector9~5_combout\ : std_logic;
SIGNAL \ALT_INV_Selector9~4_combout\ : std_logic;
SIGNAL \ALT_INV_Selector9~3_combout\ : std_logic;
SIGNAL \ALT_INV_Selector9~2_combout\ : std_logic;
SIGNAL \ALT_INV_Selector9~1_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~39_combout\ : std_logic;
SIGNAL \ALT_INV_Selector9~0_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight0~12_combout\ : std_logic;
SIGNAL \ALT_INV_Selector10~4_combout\ : std_logic;
SIGNAL \ALT_INV_Selector10~3_combout\ : std_logic;
SIGNAL \ALT_INV_Selector10~2_combout\ : std_logic;
SIGNAL \ALT_INV_Selector10~1_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~37_combout\ : std_logic;
SIGNAL \ALT_INV_Selector10~0_combout\ : std_logic;
SIGNAL \ALT_INV_Selector11~5_combout\ : std_logic;
SIGNAL \ALT_INV_Selector11~4_combout\ : std_logic;
SIGNAL \ALT_INV_Selector11~3_combout\ : std_logic;
SIGNAL \ALT_INV_Selector11~2_combout\ : std_logic;
SIGNAL \ALT_INV_Selector11~1_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~35_combout\ : std_logic;
SIGNAL \ALT_INV_Selector11~0_combout\ : std_logic;
SIGNAL \ALT_INV_vAluRes~17_combout\ : std_logic;
SIGNAL \ALT_INV_Selector12~5_combout\ : std_logic;
SIGNAL \ALT_INV_Selector12~4_combout\ : std_logic;
SIGNAL \ALT_INV_Selector12~3_combout\ : std_logic;
SIGNAL \ALT_INV_Selector12~1_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~33_combout\ : std_logic;
SIGNAL \ALT_INV_Selector12~0_combout\ : std_logic;
SIGNAL \ALT_INV_Selector13~1_combout\ : std_logic;
SIGNAL \ALT_INV_Selector13~0_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~31_combout\ : std_logic;
SIGNAL \ALT_INV_Selector14~3_combout\ : std_logic;
SIGNAL \ALT_INV_Selector14~2_combout\ : std_logic;
SIGNAL \ALT_INV_Selector14~1_combout\ : std_logic;
SIGNAL \ALT_INV_Selector14~0_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~29_combout\ : std_logic;
SIGNAL \ALT_INV_Selector15~4_combout\ : std_logic;
SIGNAL \ALT_INV_Selector15~3_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~27_combout\ : std_logic;
SIGNAL \ALT_INV_Selector15~1_combout\ : std_logic;
SIGNAL \ALT_INV_Selector15~0_combout\ : std_logic;
SIGNAL \ALT_INV_Selector16~4_combout\ : std_logic;
SIGNAL \ALT_INV_Selector16~3_combout\ : std_logic;
SIGNAL \ALT_INV_Selector16~2_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~25_combout\ : std_logic;
SIGNAL \ALT_INV_Selector17~3_combout\ : std_logic;
SIGNAL \ALT_INV_Selector17~2_combout\ : std_logic;
SIGNAL \ALT_INV_Selector17~1_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~54_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~23_combout\ : std_logic;
SIGNAL \ALT_INV_Selector18~4_combout\ : std_logic;
SIGNAL \ALT_INV_Selector18~3_combout\ : std_logic;
SIGNAL \ALT_INV_Selector18~2_combout\ : std_logic;
SIGNAL \ALT_INV_Selector18~0_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~53_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~21_combout\ : std_logic;
SIGNAL \ALT_INV_Selector19~3_combout\ : std_logic;
SIGNAL \ALT_INV_Selector19~2_combout\ : std_logic;
SIGNAL \ALT_INV_Selector19~1_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~52_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~19_combout\ : std_logic;
SIGNAL \ALT_INV_Selector20~4_combout\ : std_logic;
SIGNAL \ALT_INV_Selector20~3_combout\ : std_logic;
SIGNAL \ALT_INV_Selector20~2_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~51_combout\ : std_logic;
SIGNAL \ALT_INV_Selector20~1_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~17_combout\ : std_logic;
SIGNAL \ALT_INV_Selector21~3_combout\ : std_logic;
SIGNAL \ALT_INV_Selector21~2_combout\ : std_logic;
SIGNAL \ALT_INV_Selector21~1_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~50_combout\ : std_logic;
SIGNAL \ALT_INV_Selector21~0_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~15_combout\ : std_logic;
SIGNAL \ALT_INV_vAluRes~10_combout\ : std_logic;
SIGNAL \ALT_INV_Selector22~4_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~49_combout\ : std_logic;
SIGNAL \ALT_INV_Selector22~3_combout\ : std_logic;
SIGNAL \ALT_INV_Selector22~2_combout\ : std_logic;
SIGNAL \ALT_INV_Selector23~5_combout\ : std_logic;
SIGNAL \ALT_INV_Selector23~4_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~47_combout\ : std_logic;
SIGNAL \ALT_INV_Selector23~2_combout\ : std_logic;
SIGNAL \ALT_INV_Selector23~1_combout\ : std_logic;
SIGNAL \ALT_INV_Selector23~0_combout\ : std_logic;
SIGNAL \ALT_INV_vAluRes~8_combout\ : std_logic;
SIGNAL \ALT_INV_Selector24~3_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~46_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight0~10_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~11_combout\ : std_logic;
SIGNAL \ALT_INV_Selector24~1_combout\ : std_logic;
SIGNAL \ALT_INV_vAluRes~7_combout\ : std_logic;
SIGNAL \ALT_INV_Selector25~4_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~45_combout\ : std_logic;
SIGNAL \ALT_INV_Selector25~2_combout\ : std_logic;
SIGNAL \ALT_INV_Selector25~1_combout\ : std_logic;
SIGNAL \ALT_INV_vAluRes~6_combout\ : std_logic;
SIGNAL \ALT_INV_Selector26~3_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~44_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight0~9_combout\ : std_logic;
SIGNAL \ALT_INV_Selector26~1_combout\ : std_logic;
SIGNAL \ALT_INV_Selector26~0_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~43_combout\ : std_logic;
SIGNAL \ALT_INV_vAluRes~5_combout\ : std_logic;
SIGNAL \ALT_INV_Selector27~4_combout\ : std_logic;
SIGNAL \ALT_INV_Selector27~3_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~42_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight0~8_combout\ : std_logic;
SIGNAL \ALT_INV_Selector27~1_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~41_combout\ : std_logic;
SIGNAL \ALT_INV_vAluRes~4_combout\ : std_logic;
SIGNAL \ALT_INV_Selector28~3_combout\ : std_logic;
SIGNAL \ALT_INV_Selector28~2_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~40_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight0~6_combout\ : std_logic;
SIGNAL \ALT_INV_Selector28~0_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~39_combout\ : std_logic;
SIGNAL \ALT_INV_vAluRes~3_combout\ : std_logic;
SIGNAL \ALT_INV_Selector29~3_combout\ : std_logic;
SIGNAL \ALT_INV_Selector29~2_combout\ : std_logic;
SIGNAL \ALT_INV_Selector29~1_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~38_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~33_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight0~5_combout\ : std_logic;
SIGNAL \ALT_INV_vAluRes~2_combout\ : std_logic;
SIGNAL \ALT_INV_Selector30~3_combout\ : std_logic;
SIGNAL \ALT_INV_Selector30~2_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight0~3_combout\ : std_logic;
SIGNAL \ALT_INV_Selector30~0_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~29_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~24_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~20_combout\ : std_logic;
SIGNAL \ALT_INV_vAluRes~1_combout\ : std_logic;
SIGNAL \ALT_INV_Selector31~4_combout\ : std_logic;
SIGNAL \ALT_INV_Selector31~3_combout\ : std_logic;
SIGNAL \ALT_INV_Selector31~1_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~19_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight0~1_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~14_combout\ : std_logic;
SIGNAL \ALT_INV_vAluRes~0_combout\ : std_logic;
SIGNAL \ALT_INV_Selector32~7_combout\ : std_logic;
SIGNAL \ALT_INV_R.aluOp.ALUOpAnd~q\ : std_logic;
SIGNAL \ALT_INV_R.aluOp.ALUOpOr~q\ : std_logic;
SIGNAL \ALT_INV_R.aluOp.ALUOpSLL~q\ : std_logic;
SIGNAL \ALT_INV_R.aluOp.ALUOpSub~q\ : std_logic;
SIGNAL \ALT_INV_Selector32~2_combout\ : std_logic;
SIGNAL \ALT_INV_R.aluOp.ALUOpAdd~q\ : std_logic;
SIGNAL \ALT_INV_R.aluOp.ALUOpXor~q\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~9_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~4_combout\ : std_logic;
SIGNAL \ALT_INV_R.aluOp.ALUOpSRA~q\ : std_logic;
SIGNAL \ALT_INV_R.aluOp.ALUOpSRL~q\ : std_logic;
SIGNAL \ALT_INV_Selector32~1_combout\ : std_logic;
SIGNAL \ALT_INV_LessThan1~38_combout\ : std_logic;
SIGNAL \ALT_INV_LessThan1~37_combout\ : std_logic;
SIGNAL \ALT_INV_R.aluData2\ : std_logic_vector(31 DOWNTO 0);
SIGNAL \ALT_INV_R.aluData1\ : std_logic_vector(31 DOWNTO 2);
SIGNAL \ALT_INV_LessThan1~36_combout\ : std_logic;
SIGNAL \ALT_INV_LessThan1~35_combout\ : std_logic;
SIGNAL \ALT_INV_LessThan1~33_combout\ : std_logic;
SIGNAL \ALT_INV_LessThan1~32_combout\ : std_logic;
SIGNAL \ALT_INV_LessThan1~31_combout\ : std_logic;
SIGNAL \ALT_INV_LessThan1~27_combout\ : std_logic;
SIGNAL \ALT_INV_LessThan1~26_combout\ : std_logic;
SIGNAL \ALT_INV_LessThan1~23_combout\ : std_logic;
SIGNAL \ALT_INV_LessThan1~19_combout\ : std_logic;
SIGNAL \ALT_INV_LessThan1~17_combout\ : std_logic;
SIGNAL \ALT_INV_LessThan1~13_combout\ : std_logic;
SIGNAL \ALT_INV_LessThan1~6_combout\ : std_logic;
SIGNAL \ALT_INV_Selector32~0_combout\ : std_logic;
SIGNAL \ALT_INV_R.aluOp.ALUOpSLT~q\ : std_logic;
SIGNAL \ALT_INV_R.aluOp.ALUOpSLTU~q\ : std_logic;
SIGNAL \ALT_INV_Comb~0_combout\ : std_logic;
SIGNAL \ALT_INV_R.ctrlState.WriteReg~q\ : std_logic;
SIGNAL \ALT_INV_R.ctrlState.Wait1~q\ : std_logic;
SIGNAL \ALT_INV_vAluRes~60_combout\ : std_logic;
SIGNAL \ALT_INV_vAluRes~56_combout\ : std_logic;
SIGNAL \ALT_INV_vAluRes~52_combout\ : std_logic;
SIGNAL \ALT_INV_Selector7~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux98~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux114~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux122~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux97~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux113~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux121~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux96~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux112~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux120~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux95~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux111~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux119~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux94~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux110~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux118~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux93~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux109~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux117~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux92~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux108~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux116~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux91~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux107~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux115~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux106~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux105~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux104~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux103~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux102~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux101~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux100~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux99~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux19~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux69~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux70~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux71~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux72~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux73~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux74~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux75~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux76~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux79~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux80~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux77~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux78~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux81~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux82~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux83~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux84~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux90~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux89~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux87~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux88~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux85~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux86~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux65~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux62~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux63~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux64~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux66~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux67~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux68~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux59~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux60~26_combout\ : std_logic;
SIGNAL \ALT_INV_Mux61~26_combout\ : std_logic;
SIGNAL \ALT_INV_Add1~129_sumout\ : std_logic;
SIGNAL \ALT_INV_Add2~129_sumout\ : std_logic;
SIGNAL \ALT_INV_R.csrRead~q\ : std_logic;
SIGNAL \ALT_INV_R.memToReg~q\ : std_logic;
SIGNAL \ALT_INV_Mux61~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux61~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux61~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux60~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux60~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux60~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux59~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux59~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux59~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux68~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux68~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux68~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux67~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux67~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux67~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux66~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux66~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux66~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux64~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux64~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux64~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux63~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux63~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux63~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux62~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux62~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux62~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux65~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux65~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux65~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux86~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux86~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux86~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux85~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux85~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux85~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux88~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux88~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux88~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux87~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux87~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux87~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux89~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux89~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux89~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux90~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux90~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux90~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux84~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux84~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux84~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux83~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux83~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux83~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux82~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux82~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux82~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux81~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux81~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux81~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux78~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux78~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux78~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux77~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux77~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux77~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux80~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux80~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux80~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux79~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux79~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux79~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux76~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux76~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux76~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux75~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux75~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux75~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux74~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux74~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux74~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux73~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux73~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux73~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux72~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux72~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux72~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux71~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux71~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux71~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux70~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux70~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux70~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux69~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux69~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux69~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux99~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux99~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux99~14_combout\ : std_logic;
SIGNAL \ALT_INV_R.regWriteData\ : std_logic_vector(31 DOWNTO 0);
SIGNAL \ALT_INV_Mux100~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux100~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux100~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux101~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux101~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux101~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux102~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux102~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux102~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux103~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux103~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux103~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux104~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux104~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux104~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux105~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux105~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux105~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux106~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux106~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux106~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux115~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux115~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux115~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux107~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux107~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux107~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux91~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux91~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux91~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux116~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux116~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux116~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux108~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux108~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux108~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux92~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux92~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux92~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux117~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux117~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux117~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux109~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux109~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux109~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux93~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux93~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux93~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux118~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux118~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux118~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux110~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux110~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux110~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux94~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux94~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux94~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux119~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux119~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux119~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux111~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux111~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux111~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux95~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux95~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux95~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux120~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux120~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux120~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux112~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux112~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux112~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux96~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux96~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux96~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux121~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux121~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux121~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux113~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux113~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux113~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux97~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux97~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux97~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux122~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux122~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux122~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux114~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux114~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux114~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux98~22_combout\ : std_logic;
SIGNAL \ALT_INV_Mux98~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux98~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux61~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux61~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux61~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux60~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux60~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux60~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux59~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux59~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux59~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux68~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux68~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux68~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux67~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux67~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux67~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux66~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux66~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux66~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux64~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux64~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux64~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux63~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux63~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux63~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux62~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux62~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux62~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux65~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux65~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux65~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux86~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux86~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux86~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux85~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux85~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux85~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux88~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux88~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux88~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux87~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux87~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux87~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux89~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux89~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux89~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux90~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux90~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux90~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux84~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux84~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux84~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux83~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux83~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux83~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux82~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux82~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux82~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux81~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux81~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux81~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux78~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux78~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux78~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux77~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux77~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux77~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux80~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux80~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux80~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux79~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux79~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux79~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux76~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux76~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux76~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux75~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux75~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux75~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux74~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux74~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux74~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux73~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux73~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux73~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux72~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux72~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux72~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux71~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux71~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux71~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux70~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux70~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux70~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux69~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux69~5_combout\ : std_logic;
SIGNAL \ALT_INV_Mux69~1_combout\ : std_logic;
SIGNAL \ALT_INV_Add3~125_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~121_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~117_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~113_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~109_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~105_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~101_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~97_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~93_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~89_sumout\ : std_logic;
SIGNAL \ALT_INV_Add0~77_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~85_sumout\ : std_logic;
SIGNAL \ALT_INV_Add0~73_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~81_sumout\ : std_logic;
SIGNAL \ALT_INV_Add0~69_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~77_sumout\ : std_logic;
SIGNAL \ALT_INV_Add0~65_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~73_sumout\ : std_logic;
SIGNAL \ALT_INV_Add0~61_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~69_sumout\ : std_logic;
SIGNAL \ALT_INV_Add0~57_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~65_sumout\ : std_logic;
SIGNAL \ALT_INV_Add0~53_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~61_sumout\ : std_logic;
SIGNAL \ALT_INV_Add0~49_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~57_sumout\ : std_logic;
SIGNAL \ALT_INV_Add0~45_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~53_sumout\ : std_logic;
SIGNAL \ALT_INV_Add0~41_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~49_sumout\ : std_logic;
SIGNAL \ALT_INV_Add0~37_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~45_sumout\ : std_logic;
SIGNAL \ALT_INV_Add0~33_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~41_sumout\ : std_logic;
SIGNAL \ALT_INV_Add0~29_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~37_sumout\ : std_logic;
SIGNAL \ALT_INV_Add0~25_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~33_sumout\ : std_logic;
SIGNAL \ALT_INV_Add0~21_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~29_sumout\ : std_logic;
SIGNAL \ALT_INV_Add0~17_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~25_sumout\ : std_logic;
SIGNAL \ALT_INV_Add0~13_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~21_sumout\ : std_logic;
SIGNAL \ALT_INV_Add0~9_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~17_sumout\ : std_logic;
SIGNAL \ALT_INV_Add0~5_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~13_sumout\ : std_logic;
SIGNAL \ALT_INV_R.incPC~q\ : std_logic;
SIGNAL \ALT_INV_Add0~1_sumout\ : std_logic;
SIGNAL \ALT_INV_Add3~9_sumout\ : std_logic;
SIGNAL \ALT_INV_ShiftRight0~7_OTERM233DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][23]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][20]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][18]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][31]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][5]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][11]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][27]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][10]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][26]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][9]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][0]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][8]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][8]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][20]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][18]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][16]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][16]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][16]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][7]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][6]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][30]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][2]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][10]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][1]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][9]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][9]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][0]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][0]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][8]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_R.ctrlState.DataAccess0~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][20]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][19]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][18]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[4][18]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][17]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[5][16]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][7]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][15]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][14]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[1][29]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][12]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][28]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[2][26]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[7][26]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_RegFile[6][8]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_R.aluRes[30]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_R.aluRes[27]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_R.aluRes[4]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_R.aluRes[0]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_R.aluOp.ALUOpAnd~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_R.aluOp.ALUOpXor~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_R.aluData2[25]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_R.aluData2[13]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_R.curPC[0]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_R.curPC[31]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_R.curPC[30]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_R.curPC[21]~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[18]~1_RESYN1740_BDD1741\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[18]~1_RESYN1738_BDD1739\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[18]~1_RESYN1736_BDD1737\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[8]~1_RESYN1734_BDD1735\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[8]~1_RESYN1732_BDD1733\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[8]~1_RESYN1730_BDD1731\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[16]~0_RESYN1728_BDD1729\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[16]~0_RESYN1726_BDD1727\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[16]~0_RESYN1724_BDD1725\ : std_logic;
SIGNAL \ALT_INV_vAluRes~7_RESYN1076_RESYN1132_BDD1133\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[21]~1_RESYN1130_BDD1131\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[21]~1_RESYN1128_BDD1129\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[21]~1_RESYN1126_BDD1127\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[17]~1_RESYN1124_BDD1125\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[17]~1_RESYN1122_BDD1123\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[17]~1_RESYN1120_BDD1121\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[7]~0_RESYN1118_BDD1119\ : std_logic;
SIGNAL \ALT_INV_Selector25~6_RESYN1116_BDD1117\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[23]~2_RESYN1114_BDD1115\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[22]~2_RESYN1112_BDD1113\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[20]~2_RESYN1110_BDD1111\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[27]~2_RESYN1108_BDD1109\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[25]~2_RESYN1106_BDD1107\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[24]~3_RESYN1104_BDD1105\ : std_logic;
SIGNAL \ALT_INV_Equal3~5_RESYN1102_BDD1103\ : std_logic;
SIGNAL \ALT_INV_Equal3~5_RESYN1100_BDD1101\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[6]~0_RESYN1098_BDD1099\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[14]~1_RESYN1096_BDD1097\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[14]~1_RESYN1094_BDD1095\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[5]~0_RESYN1092_BDD1093\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[4]~0_RESYN1090_BDD1091\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[12]~1_RESYN1088_BDD1089\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[12]~1_RESYN1086_BDD1087\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[3]~0_RESYN1084_BDD1085\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[2]~0_RESYN1082_BDD1083\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[9]~1_RESYN1080_BDD1081\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[9]~1_RESYN1078_BDD1079\ : std_logic;
SIGNAL \ALT_INV_vAluRes~7_RESYN1076_BDD1077\ : std_logic;
SIGNAL \ALT_INV_vAluRes~6_RESYN1072_BDD1073\ : std_logic;
SIGNAL \ALT_INV_vAluRes~5_RESYN1070_BDD1071\ : std_logic;
SIGNAL \ALT_INV_vAluRes~4_RESYN1068_BDD1069\ : std_logic;
SIGNAL \ALT_INV_vAluRes~3_RESYN1066_BDD1067\ : std_logic;
SIGNAL \ALT_INV_vAluRes~2_RESYN1064_BDD1065\ : std_logic;
SIGNAL \ALT_INV_vAluRes~1_RESYN1062_BDD1063\ : std_logic;
SIGNAL \ALT_INV_Selector32~7_RESYN1060_BDD1061\ : std_logic;
SIGNAL \ALT_INV_Selector32~7_RESYN1058_BDD1059\ : std_logic;
SIGNAL \ALT_INV_Selector32~7_RESYN1056_BDD1057\ : std_logic;
SIGNAL \ALT_INV_Equal3~12_RESYN1054_BDD1055\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[15]~1_RESYN1048_BDD1049\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[15]~1_RESYN1046_BDD1047\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[13]~1_RESYN1044_BDD1045\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[13]~1_RESYN1042_BDD1043\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[11]~1_RESYN1040_BDD1041\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[11]~1_RESYN1038_BDD1039\ : std_logic;
SIGNAL \ALT_INV_Comb:vJumpAdr[30]~0_RESYN1036_BDD1037\ : std_logic;
SIGNAL \ALT_INV_Comb:vJumpAdr[29]~0_RESYN1034_BDD1035\ : std_logic;
SIGNAL \ALT_INV_Comb:vJumpAdr[28]~0_RESYN1032_BDD1033\ : std_logic;
SIGNAL \ALT_INV_Comb:vJumpAdr[27]~0_RESYN1030_BDD1031\ : std_logic;
SIGNAL \ALT_INV_Comb:vJumpAdr[22]~0_RESYN1028_BDD1029\ : std_logic;
SIGNAL \ALT_INV_Add2~17_OTERM727_OTERM841\ : std_logic;
SIGNAL \ALT_INV_Add2~1_OTERM735_OTERM839\ : std_logic;
SIGNAL \ALT_INV_Add2~1_OTERM735_OTERM837\ : std_logic;
SIGNAL \ALT_INV_Add2~25_OTERM723_OTERM835\ : std_logic;
SIGNAL \ALT_INV_Add2~25_OTERM723_OTERM833\ : std_logic;
SIGNAL \ALT_INV_Add2~25_OTERM723_OTERM831\ : std_logic;
SIGNAL \ALT_INV_Add2~25_OTERM723_OTERM829\ : std_logic;
SIGNAL \ALT_INV_Add2~33_OTERM719_OTERM827\ : std_logic;
SIGNAL \ALT_INV_Add2~33_OTERM719_OTERM825\ : std_logic;
SIGNAL \ALT_INV_Add2~33_OTERM719_OTERM823\ : std_logic;
SIGNAL \ALT_INV_Add2~33_OTERM719_OTERM821\ : std_logic;
SIGNAL \ALT_INV_Add2~41_OTERM715_OTERM819\ : std_logic;
SIGNAL \ALT_INV_Add2~41_OTERM715_OTERM817\ : std_logic;
SIGNAL \ALT_INV_Add2~57_OTERM707_OTERM815\ : std_logic;
SIGNAL \ALT_INV_Add2~57_OTERM707_OTERM813\ : std_logic;
SIGNAL \ALT_INV_Add2~65_OTERM703_OTERM811\ : std_logic;
SIGNAL \ALT_INV_Add2~65_OTERM703_OTERM809\ : std_logic;
SIGNAL \ALT_INV_Add2~65_OTERM703_OTERM807\ : std_logic;
SIGNAL \ALT_INV_Add2~65_OTERM703_OTERM805\ : std_logic;
SIGNAL \ALT_INV_Selector19~1_OTERM751_OTERM803\ : std_logic;
SIGNAL \ALT_INV_Selector25~3_OTERM797\ : std_logic;
SIGNAL \ALT_INV_Selector16~1_OTERM793\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~12_OTERM791\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~38_OTERM789\ : std_logic;
SIGNAL \ALT_INV_Selector1~0_OTERM771\ : std_logic;
SIGNAL \ALT_INV_Selector20~0_OTERM769\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~55_OTERM767\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~53_OTERM765\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~51_OTERM763\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~49_OTERM761\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~47_OTERM759\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~45_OTERM757\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~40_OTERM755\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~14_OTERM753\ : std_logic;
SIGNAL \ALT_INV_Selector22~0_OTERM475_OTERM749\ : std_logic;
SIGNAL \ALT_INV_Selector22~0_OTERM475_OTERM747\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~38_OTERM439_OTERM745\ : std_logic;
SIGNAL \ALT_INV_Selector15~2_OTERM741\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~26_OTERM739\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~22_OTERM737\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~36_OTERM603\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~30_OTERM601\ : std_logic;
SIGNAL \ALT_INV_Selector31~5_OTERM599\ : std_logic;
SIGNAL \ALT_INV_R.statusReg[0]_OTERM11_OTERM377_OTERM597\ : std_logic;
SIGNAL \ALT_INV_R.statusReg[0]_OTERM11_OTERM377_OTERM595\ : std_logic;
SIGNAL \ALT_INV_R.statusReg[0]_OTERM11_OTERM377_OTERM593\ : std_logic;
SIGNAL \ALT_INV_Selector31~0_NEW_REG348_OTERM569\ : std_logic;
SIGNAL \ALT_INV_R.statusReg[0]_OTERM7_OTERM491\ : std_logic;
SIGNAL \ALT_INV_R.statusReg[0]_OTERM7_OTERM489\ : std_logic;
SIGNAL \ALT_INV_R.statusReg[0]_OTERM7_OTERM487\ : std_logic;
SIGNAL \ALT_INV_R.statusReg[0]_OTERM7_OTERM485\ : std_logic;
SIGNAL \ALT_INV_R.statusReg[0]_OTERM7_OTERM483\ : std_logic;
SIGNAL \ALT_INV_R.statusReg[0]_OTERM7_OTERM481\ : std_logic;
SIGNAL \ALT_INV_Selector22~0_RTM0477_combout\ : std_logic;
SIGNAL \ALT_INV_R.statusReg[0]_OTERM9_OTERM473\ : std_logic;
SIGNAL \ALT_INV_R.statusReg[0]_OTERM9_OTERM471\ : std_logic;
SIGNAL \ALT_INV_R.statusReg[0]_OTERM9_OTERM469\ : std_logic;
SIGNAL \ALT_INV_R.statusReg[0]_OTERM9_OTERM467\ : std_logic;
SIGNAL \ALT_INV_R.statusReg[0]_OTERM9_OTERM465\ : std_logic;
SIGNAL \ALT_INV_R.statusReg[0]_OTERM9_OTERM463\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~9_OTERM461\ : std_logic;
SIGNAL \ALT_INV_Selector18~1_OTERM431\ : std_logic;
SIGNAL \ALT_INV_Selector22~1_OTERM427\ : std_logic;
SIGNAL \ALT_INV_Selector23~3_OTERM423\ : std_logic;
SIGNAL \ALT_INV_Selector24~0_OTERM419\ : std_logic;
SIGNAL \ALT_INV_Selector26~2_OTERM415\ : std_logic;
SIGNAL \ALT_INV_Selector27~2_OTERM411\ : std_logic;
SIGNAL \ALT_INV_Selector29~0_OTERM407\ : std_logic;
SIGNAL \ALT_INV_Selector30~1_OTERM403\ : std_logic;
SIGNAL \ALT_INV_Selector31~2_OTERM399\ : std_logic;
SIGNAL \ALT_INV_Selector32~4_OTERM397\ : std_logic;
SIGNAL \ALT_INV_Selector12~2_OTERM395\ : std_logic;
SIGNAL \ALT_INV_Selector16~0_OTERM393\ : std_logic;
SIGNAL \ALT_INV_Selector17~0_OTERM391\ : std_logic;
SIGNAL \ALT_INV_Selector28~1_OTERM387\ : std_logic;
SIGNAL \ALT_INV_Selector27~0_OTERM385\ : std_logic;
SIGNAL \ALT_INV_Selector31~7_OTERM383\ : std_logic;
SIGNAL \ALT_INV_Selector31~6_OTERM381\ : std_logic;
SIGNAL \ALT_INV_Selector32~3_OTERM379\ : std_logic;
SIGNAL \ALT_INV_R.statusReg[0]_OTERM11_OTERM375\ : std_logic;
SIGNAL \ALT_INV_R.statusReg[0]_OTERM11_OTERM373\ : std_logic;
SIGNAL \ALT_INV_R.statusReg[0]_OTERM11_OTERM371\ : std_logic;
SIGNAL \ALT_INV_R.statusReg[0]_OTERM11_OTERM369\ : std_logic;
SIGNAL \ALT_INV_R.statusReg[0]_OTERM11_OTERM367\ : std_logic;
SIGNAL \ALT_INV_R.aluOp.ALUOpSRA_OTERM363\ : std_logic;
SIGNAL \ALT_INV_R.aluOp.ALUOpSRL_OTERM361\ : std_logic;
SIGNAL \ALT_INV_R.aluOp.ALUOpSLL_OTERM359\ : std_logic;
SIGNAL \ALT_INV_R.aluOp.ALUOpAnd_OTERM357\ : std_logic;
SIGNAL \ALT_INV_R.aluOp.ALUOpXor_OTERM355\ : std_logic;
SIGNAL \ALT_INV_R.aluOp.ALUOpOr_OTERM353\ : std_logic;
SIGNAL \ALT_INV_Selector31~0_OTERM349\ : std_logic;
SIGNAL \ALT_INV_LessThan1~22_OTERM347\ : std_logic;
SIGNAL \ALT_INV_LessThan1~0_OTERM343\ : std_logic;
SIGNAL \ALT_INV_LessThan1~20_OTERM341\ : std_logic;
SIGNAL \ALT_INV_LessThan1~1_OTERM337\ : std_logic;
SIGNAL \ALT_INV_LessThan1~21_OTERM335\ : std_logic;
SIGNAL \ALT_INV_LessThan1~2_OTERM331\ : std_logic;
SIGNAL \ALT_INV_LessThan1~24_OTERM329\ : std_logic;
SIGNAL \ALT_INV_LessThan1~3_OTERM325\ : std_logic;
SIGNAL \ALT_INV_LessThan1~18_OTERM321\ : std_logic;
SIGNAL \ALT_INV_LessThan1~4_OTERM319\ : std_logic;
SIGNAL \ALT_INV_LessThan1~25_OTERM317\ : std_logic;
SIGNAL \ALT_INV_LessThan1~5_OTERM313\ : std_logic;
SIGNAL \ALT_INV_LessThan1~16_OTERM311\ : std_logic;
SIGNAL \ALT_INV_LessThan1~7_OTERM307\ : std_logic;
SIGNAL \ALT_INV_LessThan1~14_OTERM305\ : std_logic;
SIGNAL \ALT_INV_LessThan1~8_OTERM301\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~34_OTERM299\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~32_OTERM297\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~28_OTERM295\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~24_OTERM293\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~20_OTERM291\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~18_OTERM289\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~16_OTERM287\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~13_OTERM285\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~37_OTERM283\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~36_OTERM281\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~35_OTERM279\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~25_OTERM277\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~23_OTERM275\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~22_OTERM273\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~21_OTERM271\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~18_OTERM269\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~17_OTERM267\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~10_OTERM265\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~0_OTERM263\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~8_OTERM261\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~7_OTERM259\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~0_OTERM257\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~1_OTERM255\ : std_logic;
SIGNAL \ALT_INV_LessThan1~9_OTERM253\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~6_OTERM243\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~4_OTERM237\ : std_logic;
SIGNAL \ALT_INV_ShiftRight0~7_OTERM233\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~3_OTERM223\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~2_OTERM221\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~5_OTERM219\ : std_logic;
SIGNAL \ALT_INV_LessThan1~11_OTERM217\ : std_logic;
SIGNAL \ALT_INV_LessThan1~10_OTERM213\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~10_OTERM211\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~16_OTERM209\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~8_OTERM207\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~7_OTERM205\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~5_OTERM203\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~15_OTERM199\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~6_OTERM197\ : std_logic;
SIGNAL \ALT_INV_LessThan1~15_OTERM195\ : std_logic;
SIGNAL \ALT_INV_LessThan1~12_OTERM191\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~12_OTERM57\ : std_logic;
SIGNAL \ALT_INV_LessThan1~34_OTERM55\ : std_logic;
SIGNAL \ALT_INV_LessThan1~28_OTERM51\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~2_OTERM49\ : std_logic;
SIGNAL \ALT_INV_LessThan1~29_OTERM47\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~31_OTERM45\ : std_logic;
SIGNAL \ALT_INV_LessThan1~30_OTERM43\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~42_OTERM41\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~30_OTERM39\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~26_OTERM37\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~11_OTERM35\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~1_OTERM33\ : std_logic;
SIGNAL \ALT_INV_ShiftRight0~4_OTERM31\ : std_logic;
SIGNAL \ALT_INV_ShiftRight0~2_OTERM25\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~28_OTERM23\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~32_OTERM21\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~27_OTERM19\ : std_logic;
SIGNAL \ALT_INV_ShiftRight0~0_OTERM17\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~13_OTERM15\ : std_logic;
SIGNAL \ALT_INV_ShiftRight1~3_OTERM13\ : std_logic;
SIGNAL \ALT_INV_R.statusReg[0]_OTERM5\ : std_logic;
SIGNAL \ALT_INV_R.statusReg[0]_OTERM3\ : std_logic;
SIGNAL \ALT_INV_R.statusReg[0]_OTERM1\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[15]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[14]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[13]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[12]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[11]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[10]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[9]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[8]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[7]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[30]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[22]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[6]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[29]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[21]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[5]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[28]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[20]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[4]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[27]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[19]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[3]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[26]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[18]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[2]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[25]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[17]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[1]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[24]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[16]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[23]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[31]~input_o\ : std_logic;
SIGNAL \ALT_INV_avm_d_readdata[0]~input_o\ : std_logic;
SIGNAL \ALT_INV_Equal3~15_combout\ : std_logic;
SIGNAL \ALT_INV_Equal3~14_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[23]~3_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[23]~2_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[23]~1_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[22]~3_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[22]~2_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[22]~1_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[20]~3_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[20]~2_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[20]~1_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[27]~3_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[27]~2_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[27]~1_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[25]~3_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[25]~2_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[25]~1_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[24]~4_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[24]~3_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[24]~2_combout\ : std_logic;
SIGNAL \ALT_INV_Equal3~13_combout\ : std_logic;
SIGNAL \ALT_INV_Equal3~11_combout\ : std_logic;
SIGNAL \ALT_INV_Equal3~10_combout\ : std_logic;
SIGNAL \ALT_INV_Selector23~7_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[31]~2_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[31]~1_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[30]~2_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[30]~1_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[29]~2_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[29]~1_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[28]~2_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[28]~1_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[26]~2_combout\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[26]~1_combout\ : std_logic;
SIGNAL \ALT_INV_vAluRes~35_combout\ : std_logic;
SIGNAL \ALT_INV_vAluRes~34_combout\ : std_logic;
SIGNAL \ALT_INV_vAluRes~33_combout\ : std_logic;
SIGNAL \ALT_INV_vAluRes~32_combout\ : std_logic;
SIGNAL \ALT_INV_vAluRes~31_combout\ : std_logic;
SIGNAL \ALT_INV_Equal3~9_combout\ : std_logic;
SIGNAL \ALT_INV_Selector13~5_combout\ : std_logic;
SIGNAL \ALT_INV_Selector13~4_combout\ : std_logic;
SIGNAL \ALT_INV_Mux31~0_combout\ : std_logic;
SIGNAL \ALT_INV_Selector0~0_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~58_combout\ : std_logic;
SIGNAL \ALT_INV_ShiftLeft0~57_combout\ : std_logic;
SIGNAL \ALT_INV_Equal3~8_combout\ : std_logic;
SIGNAL \ALT_INV_Equal3~6_combout\ : std_logic;
SIGNAL \ALT_INV_Equal3~2_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][19]~q\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[19]~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][16]~q\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[24]~1_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][10]~q\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[10]~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][0]~q\ : std_logic;
SIGNAL \ALT_INV_Comb:vRegWriteData[0]~0_combout\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[26][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[24][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[27][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[25][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[18][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[16][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[19][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[17][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[10][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[8][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[11][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[9][24]~q\ : std_logic;
SIGNAL \ALT_INV_R.regWriteEn~1_combout\ : std_logic;
SIGNAL \ALT_INV_R.regWriteEn~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR~15_combout\ : std_logic;
SIGNAL \ALT_INV_Mux50~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux34~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux11~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR~10_combout\ : std_logic;
SIGNAL \ALT_INV_Mux44~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux58~0_combout\ : std_logic;
SIGNAL \ALT_INV_R.statusReg\ : std_logic_vector(2 DOWNTO 1);
SIGNAL \ALT_INV_R.ctrlState.CheckJump~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][23]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][22]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][21]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][20]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][19]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][18]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][17]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][16]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][7]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][15]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][31]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][6]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][14]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][30]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][5]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][13]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][29]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][4]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][12]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][28]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][3]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][11]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][27]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][2]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][10]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][26]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][1]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][9]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][25]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][0]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][8]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[30][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[28][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[31][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[29][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[22][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[20][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[23][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[21][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[14][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[12][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[15][24]~q\ : std_logic;
SIGNAL \ALT_INV_RegFile[13][24]~q\ : std_logic;
SIGNAL \ALT_INV_R.regWriteEn~q\ : std_logic;
SIGNAL \ALT_INV_Selector23~6_combout\ : std_logic;
SIGNAL \ALT_INV_Selector25~6_combout\ : std_logic;
SIGNAL \ALT_INV_Mux21~2_combout\ : std_logic;
SIGNAL \ALT_INV_Mux21~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux22~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux22~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux24~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux24~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux18~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux17~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux17~0_combout\ : std_logic;
SIGNAL \ALT_INV_Comb~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux0~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux23~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux23~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux26~2_combout\ : std_logic;
SIGNAL \ALT_INV_Mux26~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux25~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux25~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux21~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux125~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux225~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux61~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux61~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux124~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux224~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux60~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux60~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR.aluData2[31]~29_combout\ : std_logic;
SIGNAL \ALT_INV_Mux123~3_combout\ : std_logic;
SIGNAL \ALT_INV_Mux223~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux59~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux59~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux132~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux232~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux68~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux68~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux131~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux231~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux67~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux67~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux130~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux230~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux66~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux66~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR.aluData2[26]~25_combout\ : std_logic;
SIGNAL \ALT_INV_Mux128~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux228~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux64~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux64~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR.aluData2[27]~24_combout\ : std_logic;
SIGNAL \ALT_INV_Mux127~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux227~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux63~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux63~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR.aluData2[28]~23_combout\ : std_logic;
SIGNAL \ALT_INV_Mux126~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux226~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux62~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux62~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux129~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux229~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux65~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux65~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux250~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux86~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux86~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR.aluData2[5]~21_combout\ : std_logic;
SIGNAL \ALT_INV_Mux149~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux249~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux85~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux85~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR.aluData2[4]~20_combout\ : std_logic;
SIGNAL \ALT_INV_Mux150~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux252~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux88~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux88~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux251~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux87~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux87~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR.aluData2[2]~19_combout\ : std_logic;
SIGNAL \ALT_INV_Mux152~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR.aluData2[3]~18_combout\ : std_logic;
SIGNAL \ALT_INV_Mux151~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux253~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux89~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux89~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR.aluData2[1]~17_combout\ : std_logic;
SIGNAL \ALT_INV_Mux153~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR.aluData2[0]~16_combout\ : std_logic;
SIGNAL \ALT_INV_Mux154~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux254~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux90~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux90~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR.aluData2[6]~15_combout\ : std_logic;
SIGNAL \ALT_INV_Mux148~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux248~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux84~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux84~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR.aluData2[7]~14_combout\ : std_logic;
SIGNAL \ALT_INV_Mux147~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux247~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux83~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux83~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR.aluData2[8]~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux146~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux246~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux82~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux82~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR.aluData2[9]~12_combout\ : std_logic;
SIGNAL \ALT_INV_Mux145~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux245~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux81~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux81~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR.aluData2[12]~11_combout\ : std_logic;
SIGNAL \ALT_INV_Mux142~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux242~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux78~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux78~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR.aluData2[13]~10_combout\ : std_logic;
SIGNAL \ALT_INV_Mux141~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux241~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux77~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux77~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR.aluData2[10]~9_combout\ : std_logic;
SIGNAL \ALT_INV_Mux144~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux244~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux80~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux80~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR.aluData2[11]~8_combout\ : std_logic;
SIGNAL \ALT_INV_Mux143~1_combout\ : std_logic;
SIGNAL \ALT_INV_Mux143~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux243~0_combout\ : std_logic;
SIGNAL \ALT_INV_Mux79~13_combout\ : std_logic;
SIGNAL \ALT_INV_Mux79~0_combout\ : std_logic;
SIGNAL \ALT_INV_NxR.aluData2[14]~7_combout\ : std_logic;
SIGNAL \ALT_INV_Mux140~0_combout\ : std_logic;

BEGIN

ww_csi_clk <= csi_clk;
ww_rsi_reset_n <= rsi_reset_n;
avm_i_address <= ww_avm_i_address;
avm_i_read <= ww_avm_i_read;
ww_avm_i_readdata <= avm_i_readdata;
ww_avm_i_waitrequest <= avm_i_waitrequest;
avm_d_address <= ww_avm_d_address;
avm_d_byteenable <= ww_avm_d_byteenable;
avm_d_write <= ww_avm_d_write;
avm_d_writedata <= ww_avm_d_writedata;
avm_d_read <= ww_avm_d_read;
ww_avm_d_readdata <= avm_d_readdata;
ww_avm_d_waitrequest <= avm_d_waitrequest;
ww_devoe <= devoe;
ww_devclrn <= devclrn;
ww_devpor <= devpor;
\ALT_INV_Add3~5_sumout\ <= NOT \Add3~5_sumout\;
\ALT_INV_R.jumpToAdr~q\ <= NOT \R.jumpToAdr~q\;
\ALT_INV_Add3~1_sumout\ <= NOT \Add3~1_sumout\;
\ALT_INV_Mux99~9_combout\ <= NOT \Mux99~9_combout\;
\ALT_INV_Mux99~5_combout\ <= NOT \Mux99~5_combout\;
\ALT_INV_Mux99~1_combout\ <= NOT \Mux99~1_combout\;
\ALT_INV_Mux100~9_combout\ <= NOT \Mux100~9_combout\;
\ALT_INV_Mux100~5_combout\ <= NOT \Mux100~5_combout\;
\ALT_INV_Mux100~1_combout\ <= NOT \Mux100~1_combout\;
\ALT_INV_Mux101~9_combout\ <= NOT \Mux101~9_combout\;
\ALT_INV_Mux101~5_combout\ <= NOT \Mux101~5_combout\;
\ALT_INV_Mux101~1_combout\ <= NOT \Mux101~1_combout\;
\ALT_INV_Mux102~9_combout\ <= NOT \Mux102~9_combout\;
\ALT_INV_Mux102~5_combout\ <= NOT \Mux102~5_combout\;
\ALT_INV_Mux102~1_combout\ <= NOT \Mux102~1_combout\;
\ALT_INV_Mux103~9_combout\ <= NOT \Mux103~9_combout\;
\ALT_INV_Mux103~5_combout\ <= NOT \Mux103~5_combout\;
\ALT_INV_Mux103~1_combout\ <= NOT \Mux103~1_combout\;
\ALT_INV_Mux104~9_combout\ <= NOT \Mux104~9_combout\;
\ALT_INV_Mux104~5_combout\ <= NOT \Mux104~5_combout\;
\ALT_INV_Mux104~1_combout\ <= NOT \Mux104~1_combout\;
\ALT_INV_Mux105~9_combout\ <= NOT \Mux105~9_combout\;
\ALT_INV_Mux105~5_combout\ <= NOT \Mux105~5_combout\;
\ALT_INV_Mux105~1_combout\ <= NOT \Mux105~1_combout\;
\ALT_INV_Mux106~9_combout\ <= NOT \Mux106~9_combout\;
\ALT_INV_Mux106~5_combout\ <= NOT \Mux106~5_combout\;
\ALT_INV_Mux106~1_combout\ <= NOT \Mux106~1_combout\;
\ALT_INV_Mux115~9_combout\ <= NOT \Mux115~9_combout\;
\ALT_INV_Mux115~5_combout\ <= NOT \Mux115~5_combout\;
\ALT_INV_Mux115~1_combout\ <= NOT \Mux115~1_combout\;
\ALT_INV_Mux107~9_combout\ <= NOT \Mux107~9_combout\;
\ALT_INV_Mux107~5_combout\ <= NOT \Mux107~5_combout\;
\ALT_INV_Mux107~1_combout\ <= NOT \Mux107~1_combout\;
\ALT_INV_Mux91~9_combout\ <= NOT \Mux91~9_combout\;
\ALT_INV_Mux91~5_combout\ <= NOT \Mux91~5_combout\;
\ALT_INV_Mux91~1_combout\ <= NOT \Mux91~1_combout\;
\ALT_INV_Mux116~9_combout\ <= NOT \Mux116~9_combout\;
\ALT_INV_Mux116~5_combout\ <= NOT \Mux116~5_combout\;
\ALT_INV_Mux116~1_combout\ <= NOT \Mux116~1_combout\;
\ALT_INV_Mux108~9_combout\ <= NOT \Mux108~9_combout\;
\ALT_INV_Mux108~5_combout\ <= NOT \Mux108~5_combout\;
\ALT_INV_Mux108~1_combout\ <= NOT \Mux108~1_combout\;
\ALT_INV_Mux92~9_combout\ <= NOT \Mux92~9_combout\;
\ALT_INV_Mux92~5_combout\ <= NOT \Mux92~5_combout\;
\ALT_INV_Mux92~1_combout\ <= NOT \Mux92~1_combout\;
\ALT_INV_Mux117~9_combout\ <= NOT \Mux117~9_combout\;
\ALT_INV_Mux117~5_combout\ <= NOT \Mux117~5_combout\;
\ALT_INV_Mux117~1_combout\ <= NOT \Mux117~1_combout\;
\ALT_INV_Mux109~9_combout\ <= NOT \Mux109~9_combout\;
\ALT_INV_Mux109~5_combout\ <= NOT \Mux109~5_combout\;
\ALT_INV_Mux109~1_combout\ <= NOT \Mux109~1_combout\;
\ALT_INV_Mux93~9_combout\ <= NOT \Mux93~9_combout\;
\ALT_INV_Mux93~5_combout\ <= NOT \Mux93~5_combout\;
\ALT_INV_Mux93~1_combout\ <= NOT \Mux93~1_combout\;
\ALT_INV_Mux118~9_combout\ <= NOT \Mux118~9_combout\;
\ALT_INV_Mux118~5_combout\ <= NOT \Mux118~5_combout\;
\ALT_INV_Mux118~1_combout\ <= NOT \Mux118~1_combout\;
\ALT_INV_Mux110~9_combout\ <= NOT \Mux110~9_combout\;
\ALT_INV_Mux110~5_combout\ <= NOT \Mux110~5_combout\;
\ALT_INV_Mux110~1_combout\ <= NOT \Mux110~1_combout\;
\ALT_INV_Mux94~9_combout\ <= NOT \Mux94~9_combout\;
\ALT_INV_Mux94~5_combout\ <= NOT \Mux94~5_combout\;
\ALT_INV_Mux94~1_combout\ <= NOT \Mux94~1_combout\;
\ALT_INV_Mux119~9_combout\ <= NOT \Mux119~9_combout\;
\ALT_INV_Mux119~5_combout\ <= NOT \Mux119~5_combout\;
\ALT_INV_Mux119~1_combout\ <= NOT \Mux119~1_combout\;
\ALT_INV_Mux111~9_combout\ <= NOT \Mux111~9_combout\;
\ALT_INV_Mux111~5_combout\ <= NOT \Mux111~5_combout\;
\ALT_INV_Mux111~1_combout\ <= NOT \Mux111~1_combout\;
\ALT_INV_Mux95~9_combout\ <= NOT \Mux95~9_combout\;
\ALT_INV_Mux95~5_combout\ <= NOT \Mux95~5_combout\;
\ALT_INV_Mux95~1_combout\ <= NOT \Mux95~1_combout\;
\ALT_INV_Mux120~9_combout\ <= NOT \Mux120~9_combout\;
\ALT_INV_Mux120~5_combout\ <= NOT \Mux120~5_combout\;
\ALT_INV_Mux120~1_combout\ <= NOT \Mux120~1_combout\;
\ALT_INV_Mux112~9_combout\ <= NOT \Mux112~9_combout\;
\ALT_INV_Mux112~5_combout\ <= NOT \Mux112~5_combout\;
\ALT_INV_Mux112~1_combout\ <= NOT \Mux112~1_combout\;
\ALT_INV_Mux96~9_combout\ <= NOT \Mux96~9_combout\;
\ALT_INV_Mux96~5_combout\ <= NOT \Mux96~5_combout\;
\ALT_INV_Mux96~1_combout\ <= NOT \Mux96~1_combout\;
\ALT_INV_Mux121~9_combout\ <= NOT \Mux121~9_combout\;
\ALT_INV_Mux121~5_combout\ <= NOT \Mux121~5_combout\;
\ALT_INV_Mux121~1_combout\ <= NOT \Mux121~1_combout\;
\ALT_INV_Mux113~9_combout\ <= NOT \Mux113~9_combout\;
\ALT_INV_Mux113~5_combout\ <= NOT \Mux113~5_combout\;
\ALT_INV_Mux113~1_combout\ <= NOT \Mux113~1_combout\;
\ALT_INV_Mux97~9_combout\ <= NOT \Mux97~9_combout\;
\ALT_INV_Mux97~5_combout\ <= NOT \Mux97~5_combout\;
\ALT_INV_Mux97~1_combout\ <= NOT \Mux97~1_combout\;
\ALT_INV_Mux122~9_combout\ <= NOT \Mux122~9_combout\;
\ALT_INV_Mux122~5_combout\ <= NOT \Mux122~5_combout\;
\ALT_INV_Mux122~1_combout\ <= NOT \Mux122~1_combout\;
\ALT_INV_Mux114~9_combout\ <= NOT \Mux114~9_combout\;
\ALT_INV_Mux114~5_combout\ <= NOT \Mux114~5_combout\;
\ALT_INV_Mux114~1_combout\ <= NOT \Mux114~1_combout\;
\ALT_INV_Mux98~9_combout\ <= NOT \Mux98~9_combout\;
\ALT_INV_Mux98~5_combout\ <= NOT \Mux98~5_combout\;
\ALT_INV_Mux98~1_combout\ <= NOT \Mux98~1_combout\;
\ALT_INV_Add1~125_sumout\ <= NOT \Add1~125_sumout\;
\ALT_INV_Add2~125_sumout\ <= NOT \Add2~125_sumout\;
\ALT_INV_Add1~121_sumout\ <= NOT \Add1~121_sumout\;
\ALT_INV_Add2~121_sumout\ <= NOT \Add2~121_sumout\;
\ALT_INV_Add1~117_sumout\ <= NOT \Add1~117_sumout\;
\ALT_INV_Add2~117_sumout\ <= NOT \Add2~117_sumout\;
\ALT_INV_Add1~113_sumout\ <= NOT \Add1~113_sumout\;
\ALT_INV_Add2~113_sumout\ <= NOT \Add2~113_sumout\;
\ALT_INV_Add1~109_sumout\ <= NOT \Add1~109_sumout\;
\ALT_INV_Add2~109_sumout\ <= NOT \Add2~109_sumout\;
\ALT_INV_Add1~105_sumout\ <= NOT \Add1~105_sumout\;
\ALT_INV_Add2~105_sumout\ <= NOT \Add2~105_sumout\;
\ALT_INV_Add1~101_sumout\ <= NOT \Add1~101_sumout\;
\ALT_INV_Add2~101_sumout\ <= NOT \Add2~101_sumout\;
\ALT_INV_Add1~97_sumout\ <= NOT \Add1~97_sumout\;
\ALT_INV_Add2~97_sumout\ <= NOT \Add2~97_sumout\;
\ALT_INV_Add1~93_sumout\ <= NOT \Add1~93_sumout\;
\ALT_INV_Add2~93_sumout\ <= NOT \Add2~93_sumout\;
\ALT_INV_Add1~89_sumout\ <= NOT \Add1~89_sumout\;
\ALT_INV_Add2~89_sumout\ <= NOT \Add2~89_sumout\;
\ALT_INV_Add1~85_sumout\ <= NOT \Add1~85_sumout\;
\ALT_INV_Add2~85_sumout\ <= NOT \Add2~85_sumout\;
\ALT_INV_Add1~81_sumout\ <= NOT \Add1~81_sumout\;
\ALT_INV_Add2~81_sumout\ <= NOT \Add2~81_sumout\;
\ALT_INV_Add1~77_sumout\ <= NOT \Add1~77_sumout\;
\ALT_INV_Add2~77_sumout\ <= NOT \Add2~77_sumout\;
\ALT_INV_Add1~73_sumout\ <= NOT \Add1~73_sumout\;
\ALT_INV_Add2~73_sumout\ <= NOT \Add2~73_sumout\;
\ALT_INV_Add1~69_sumout\ <= NOT \Add1~69_sumout\;
\ALT_INV_Add2~69_sumout\ <= NOT \Add2~69_sumout\;
\ALT_INV_Add1~65_sumout\ <= NOT \Add1~65_sumout\;
\ALT_INV_Add2~65_sumout\ <= NOT \Add2~65_sumout\;
\ALT_INV_Add1~61_sumout\ <= NOT \Add1~61_sumout\;
\ALT_INV_Add2~61_sumout\ <= NOT \Add2~61_sumout\;
\ALT_INV_Add1~57_sumout\ <= NOT \Add1~57_sumout\;
\ALT_INV_Add2~57_sumout\ <= NOT \Add2~57_sumout\;
\ALT_INV_Add1~53_sumout\ <= NOT \Add1~53_sumout\;
\ALT_INV_Add2~53_sumout\ <= NOT \Add2~53_sumout\;
\ALT_INV_Add1~49_sumout\ <= NOT \Add1~49_sumout\;
\ALT_INV_Add2~49_sumout\ <= NOT \Add2~49_sumout\;
\ALT_INV_Add1~45_sumout\ <= NOT \Add1~45_sumout\;
\ALT_INV_Add2~45_sumout\ <= NOT \Add2~45_sumout\;
\ALT_INV_Add1~41_sumout\ <= NOT \Add1~41_sumout\;
\ALT_INV_Add2~41_sumout\ <= NOT \Add2~41_sumout\;
\ALT_INV_Add1~37_sumout\ <= NOT \Add1~37_sumout\;
\ALT_INV_Add2~37_sumout\ <= NOT \Add2~37_sumout\;
\ALT_INV_Add1~33_sumout\ <= NOT \Add1~33_sumout\;
\ALT_INV_Add2~33_sumout\ <= NOT \Add2~33_sumout\;
\ALT_INV_Add1~29_sumout\ <= NOT \Add1~29_sumout\;
\ALT_INV_Add2~29_sumout\ <= NOT \Add2~29_sumout\;
\ALT_INV_Add1~25_sumout\ <= NOT \Add1~25_sumout\;
\ALT_INV_Add2~25_sumout\ <= NOT \Add2~25_sumout\;
\ALT_INV_Add1~21_sumout\ <= NOT \Add1~21_sumout\;
\ALT_INV_Add2~21_sumout\ <= NOT \Add2~21_sumout\;
\ALT_INV_Add1~17_sumout\ <= NOT \Add1~17_sumout\;
\ALT_INV_Add2~17_sumout\ <= NOT \Add2~17_sumout\;
\ALT_INV_Add1~13_sumout\ <= NOT \Add1~13_sumout\;
\ALT_INV_Add2~13_sumout\ <= NOT \Add2~13_sumout\;
\ALT_INV_Add2~9_sumout\ <= NOT \Add2~9_sumout\;
\ALT_INV_Add1~9_sumout\ <= NOT \Add1~9_sumout\;
\ALT_INV_Add1~5_sumout\ <= NOT \Add1~5_sumout\;
\ALT_INV_Add2~5_sumout\ <= NOT \Add2~5_sumout\;
\ALT_INV_Add2~1_sumout\ <= NOT \Add2~1_sumout\;
\ALT_INV_R.aluCalc~q\ <= NOT \R.aluCalc~q\;
\ALT_INV_R.curPC\(31) <= NOT \R.curPC\(31);
\ALT_INV_R.curPC\(30) <= NOT \R.curPC\(30);
\ALT_INV_R.curPC\(29) <= NOT \R.curPC\(29);
\ALT_INV_R.curPC\(28) <= NOT \R.curPC\(28);
\ALT_INV_R.curPC\(27) <= NOT \R.curPC\(27);
\ALT_INV_R.curPC\(26) <= NOT \R.curPC\(26);
\ALT_INV_R.curPC\(25) <= NOT \R.curPC\(25);
\ALT_INV_R.curPC\(24) <= NOT \R.curPC\(24);
\ALT_INV_R.curPC\(23) <= NOT \R.curPC\(23);
\ALT_INV_R.curPC\(22) <= NOT \R.curPC\(22);
\ALT_INV_R.curPC\(21) <= NOT \R.curPC\(21);
\ALT_INV_R.curPC\(20) <= NOT \R.curPC\(20);
\ALT_INV_R.curPC\(19) <= NOT \R.curPC\(19);
\ALT_INV_R.curPC\(18) <= NOT \R.curPC\(18);
\ALT_INV_R.curPC\(17) <= NOT \R.curPC\(17);
\ALT_INV_R.curPC\(16) <= NOT \R.curPC\(16);
\ALT_INV_R.curPC\(15) <= NOT \R.curPC\(15);
\ALT_INV_R.curPC\(14) <= NOT \R.curPC\(14);
\ALT_INV_R.curPC\(13) <= NOT \R.curPC\(13);
\ALT_INV_R.curPC\(12) <= NOT \R.curPC\(12);
\ALT_INV_R.curPC\(11) <= NOT \R.curPC\(11);
\ALT_INV_R.curPC\(10) <= NOT \R.curPC\(10);
\ALT_INV_R.curPC\(9) <= NOT \R.curPC\(9);
\ALT_INV_R.curPC\(8) <= NOT \R.curPC\(8);
\ALT_INV_R.curPC\(7) <= NOT \R.curPC\(7);
\ALT_INV_R.curPC\(6) <= NOT \R.curPC\(6);
\ALT_INV_R.curPC\(5) <= NOT \R.curPC\(5);
\ALT_INV_R.curPC\(4) <= NOT \R.curPC\(4);
\ALT_INV_R.curPC\(3) <= NOT \R.curPC\(3);
\ALT_INV_R.curPC\(2) <= NOT \R.curPC\(2);
\ALT_INV_Mux240~0_combout\ <= NOT \Mux240~0_combout\;
\ALT_INV_Mux76~13_combout\ <= NOT \Mux76~13_combout\;
\ALT_INV_Mux76~0_combout\ <= NOT \Mux76~0_combout\;
\ALT_INV_NxR.aluData2[15]~6_combout\ <= NOT \NxR.aluData2[15]~6_combout\;
\ALT_INV_Mux139~0_combout\ <= NOT \Mux139~0_combout\;
\ALT_INV_Mux239~0_combout\ <= NOT \Mux239~0_combout\;
\ALT_INV_Mux75~13_combout\ <= NOT \Mux75~13_combout\;
\ALT_INV_Mux75~0_combout\ <= NOT \Mux75~0_combout\;
\ALT_INV_NxR.aluData2[16]~5_combout\ <= NOT \NxR.aluData2[16]~5_combout\;
\ALT_INV_Mux138~0_combout\ <= NOT \Mux138~0_combout\;
\ALT_INV_Mux238~0_combout\ <= NOT \Mux238~0_combout\;
\ALT_INV_Mux74~13_combout\ <= NOT \Mux74~13_combout\;
\ALT_INV_Mux74~0_combout\ <= NOT \Mux74~0_combout\;
\ALT_INV_NxR.aluData2[17]~4_combout\ <= NOT \NxR.aluData2[17]~4_combout\;
\ALT_INV_Mux137~0_combout\ <= NOT \Mux137~0_combout\;
\ALT_INV_Mux237~0_combout\ <= NOT \Mux237~0_combout\;
\ALT_INV_Mux73~13_combout\ <= NOT \Mux73~13_combout\;
\ALT_INV_Mux73~0_combout\ <= NOT \Mux73~0_combout\;
\ALT_INV_NxR.aluData2[18]~3_combout\ <= NOT \NxR.aluData2[18]~3_combout\;
\ALT_INV_Mux136~0_combout\ <= NOT \Mux136~0_combout\;
\ALT_INV_Mux236~0_combout\ <= NOT \Mux236~0_combout\;
\ALT_INV_Mux72~13_combout\ <= NOT \Mux72~13_combout\;
\ALT_INV_Mux72~0_combout\ <= NOT \Mux72~0_combout\;
\ALT_INV_NxR.aluData2[19]~2_combout\ <= NOT \NxR.aluData2[19]~2_combout\;
\ALT_INV_Mux135~0_combout\ <= NOT \Mux135~0_combout\;
\ALT_INV_Mux123~2_combout\ <= NOT \Mux123~2_combout\;
\ALT_INV_Mux149~0_combout\ <= NOT \Mux149~0_combout\;
\ALT_INV_Mux235~0_combout\ <= NOT \Mux235~0_combout\;
\ALT_INV_Mux71~13_combout\ <= NOT \Mux71~13_combout\;
\ALT_INV_Mux71~0_combout\ <= NOT \Mux71~0_combout\;
\ALT_INV_NxR.aluData2[20]~1_combout\ <= NOT \NxR.aluData2[20]~1_combout\;
\ALT_INV_Mux134~0_combout\ <= NOT \Mux134~0_combout\;
\ALT_INV_Mux234~0_combout\ <= NOT \Mux234~0_combout\;
\ALT_INV_Mux70~13_combout\ <= NOT \Mux70~13_combout\;
\ALT_INV_Mux70~0_combout\ <= NOT \Mux70~0_combout\;
\ALT_INV_NxR.aluData2[21]~0_combout\ <= NOT \NxR.aluData2[21]~0_combout\;
\ALT_INV_vAluSrc2~1_combout\ <= NOT \vAluSrc2~1_combout\;
\ALT_INV_Mux133~0_combout\ <= NOT \Mux133~0_combout\;
\ALT_INV_Mux123~1_combout\ <= NOT \Mux123~1_combout\;
\ALT_INV_Mux124~0_combout\ <= NOT \Mux124~0_combout\;
\ALT_INV_Mux233~0_combout\ <= NOT \Mux233~0_combout\;
\ALT_INV_Mux69~13_combout\ <= NOT \Mux69~13_combout\;
\ALT_INV_R.curInst\(19) <= NOT \R.curInst\(19);
\ALT_INV_R.curInst\(18) <= NOT \R.curInst\(18);
\ALT_INV_Mux69~0_combout\ <= NOT \Mux69~0_combout\;
\ALT_INV_R.curInst\(16) <= NOT \R.curInst\(16);
\ALT_INV_R.curInst\(15) <= NOT \R.curInst\(15);
\ALT_INV_R.curInst\(17) <= NOT \R.curInst\(17);
\ALT_INV_vAluSrc1~2_combout\ <= NOT \vAluSrc1~2_combout\;
\ALT_INV_vAluSrc1~1_combout\ <= NOT \vAluSrc1~1_combout\;
\ALT_INV_vAluSrc2~0_combout\ <= NOT \vAluSrc2~0_combout\;
\ALT_INV_Mux20~1_combout\ <= NOT \Mux20~1_combout\;
\ALT_INV_Mux20~0_combout\ <= NOT \Mux20~0_combout\;
\ALT_INV_Mux26~0_combout\ <= NOT \Mux26~0_combout\;
\ALT_INV_R.ctrlState.Fetch~q\ <= NOT \R.ctrlState.Fetch~q\;
\ALT_INV_Mux12~0_combout\ <= NOT \Mux12~0_combout\;
\ALT_INV_NxR~4_combout\ <= NOT \NxR~4_combout\;
\ALT_INV_Mux154~0_combout\ <= NOT \Mux154~0_combout\;
\ALT_INV_R.ctrlState.ReadReg~q\ <= NOT \R.ctrlState.ReadReg~q\;
\ALT_INV_NxR~2_combout\ <= NOT \NxR~2_combout\;
\ALT_INV_vAluSrc1~0_combout\ <= NOT \vAluSrc1~0_combout\;
\ALT_INV_Mux123~0_combout\ <= NOT \Mux123~0_combout\;
\ALT_INV_Mux53~2_combout\ <= NOT \Mux53~2_combout\;
\ALT_INV_R.ctrlState.DataAccess1~q\ <= NOT \R.ctrlState.DataAccess1~q\;
\ALT_INV_NxR~0_combout\ <= NOT \NxR~0_combout\;
\ALT_INV_Equal2~2_combout\ <= NOT \Equal2~2_combout\;
\ALT_INV_Equal2~1_combout\ <= NOT \Equal2~1_combout\;
\ALT_INV_R.curInst\(25) <= NOT \R.curInst\(25);
\ALT_INV_Equal2~0_combout\ <= NOT \Equal2~0_combout\;
\ALT_INV_R.curInst\(31) <= NOT \R.curInst\(31);
\ALT_INV_R.curInst\(30) <= NOT \R.curInst\(30);
\ALT_INV_R.curInst\(29) <= NOT \R.curInst\(29);
\ALT_INV_R.curInst\(28) <= NOT \R.curInst\(28);
\ALT_INV_R.curInst\(27) <= NOT \R.curInst\(27);
\ALT_INV_R.curInst\(26) <= NOT \R.curInst\(26);
\ALT_INV_R.ctrlState.Trap~q\ <= NOT \R.ctrlState.Trap~q\;
\ALT_INV_R.ctrlState.Wait0~q\ <= NOT \R.ctrlState.Wait0~q\;
\ALT_INV_Mux53~1_combout\ <= NOT \Mux53~1_combout\;
\ALT_INV_Mux53~0_combout\ <= NOT \Mux53~0_combout\;
\ALT_INV_R.ctrlState.DataAccess0~q\ <= NOT \R.ctrlState.DataAccess0~q\;
\ALT_INV_R.ctrlState.Calc~q\ <= NOT \R.ctrlState.Calc~q\;
\ALT_INV_Mux18~0_combout\ <= NOT \Mux18~0_combout\;
\ALT_INV_vAluRes~30_combout\ <= NOT \vAluRes~30_combout\;
\ALT_INV_vAluRes~29_combout\ <= NOT \vAluRes~29_combout\;
\ALT_INV_vAluRes~28_combout\ <= NOT \vAluRes~28_combout\;
\ALT_INV_vAluRes~27_combout\ <= NOT \vAluRes~27_combout\;
\ALT_INV_vAluRes~26_combout\ <= NOT \vAluRes~26_combout\;
\ALT_INV_vAluRes~25_combout\ <= NOT \vAluRes~25_combout\;
\ALT_INV_Selector7~4_combout\ <= NOT \Selector7~4_combout\;
\ALT_INV_Selector13~2_combout\ <= NOT \Selector13~2_combout\;
\ALT_INV_Selector14~4_combout\ <= NOT \Selector14~4_combout\;
\ALT_INV_Selector15~5_combout\ <= NOT \Selector15~5_combout\;
\ALT_INV_Selector16~5_combout\ <= NOT \Selector16~5_combout\;
\ALT_INV_Equal4~2_combout\ <= NOT \Equal4~2_combout\;
\ALT_INV_Equal4~1_combout\ <= NOT \Equal4~1_combout\;
\ALT_INV_R.curInst\(0) <= NOT \R.curInst\(0);
\ALT_INV_R.curInst\(1) <= NOT \R.curInst\(1);
\ALT_INV_Equal4~0_combout\ <= NOT \Equal4~0_combout\;
\ALT_INV_R.curInst\(2) <= NOT \R.curInst\(2);
\ALT_INV_R.curInst\(6) <= NOT \R.curInst\(6);
\ALT_INV_R.curInst\(4) <= NOT \R.curInst\(4);
\ALT_INV_R.curInst\(5) <= NOT \R.curInst\(5);
\ALT_INV_R.curInst\(3) <= NOT \R.curInst\(3);
\ALT_INV_Mux99~13_combout\ <= NOT \Mux99~13_combout\;
\ALT_INV_RegFile[3][23]~q\ <= NOT \RegFile[3][23]~q\;
\ALT_INV_RegFile[1][23]~q\ <= NOT \RegFile[1][23]~q\;
\ALT_INV_RegFile[2][23]~q\ <= NOT \RegFile[2][23]~q\;
\ALT_INV_Mux99~0_combout\ <= NOT \Mux99~0_combout\;
\ALT_INV_RegFile[7][23]~q\ <= NOT \RegFile[7][23]~q\;
\ALT_INV_RegFile[6][23]~q\ <= NOT \RegFile[6][23]~q\;
\ALT_INV_RegFile[5][23]~q\ <= NOT \RegFile[5][23]~q\;
\ALT_INV_RegFile[4][23]~q\ <= NOT \RegFile[4][23]~q\;
\ALT_INV_Mux100~13_combout\ <= NOT \Mux100~13_combout\;
\ALT_INV_RegFile[3][22]~q\ <= NOT \RegFile[3][22]~q\;
\ALT_INV_RegFile[1][22]~q\ <= NOT \RegFile[1][22]~q\;
\ALT_INV_RegFile[2][22]~q\ <= NOT \RegFile[2][22]~q\;
\ALT_INV_Mux100~0_combout\ <= NOT \Mux100~0_combout\;
\ALT_INV_RegFile[7][22]~q\ <= NOT \RegFile[7][22]~q\;
\ALT_INV_RegFile[6][22]~q\ <= NOT \RegFile[6][22]~q\;
\ALT_INV_RegFile[5][22]~q\ <= NOT \RegFile[5][22]~q\;
\ALT_INV_RegFile[4][22]~q\ <= NOT \RegFile[4][22]~q\;
\ALT_INV_Mux101~13_combout\ <= NOT \Mux101~13_combout\;
\ALT_INV_RegFile[3][21]~q\ <= NOT \RegFile[3][21]~q\;
\ALT_INV_RegFile[1][21]~q\ <= NOT \RegFile[1][21]~q\;
\ALT_INV_RegFile[2][21]~q\ <= NOT \RegFile[2][21]~q\;
\ALT_INV_Mux101~0_combout\ <= NOT \Mux101~0_combout\;
\ALT_INV_RegFile[7][21]~q\ <= NOT \RegFile[7][21]~q\;
\ALT_INV_RegFile[6][21]~q\ <= NOT \RegFile[6][21]~q\;
\ALT_INV_RegFile[5][21]~q\ <= NOT \RegFile[5][21]~q\;
\ALT_INV_RegFile[4][21]~q\ <= NOT \RegFile[4][21]~q\;
\ALT_INV_Mux102~13_combout\ <= NOT \Mux102~13_combout\;
\ALT_INV_RegFile[3][20]~q\ <= NOT \RegFile[3][20]~q\;
\ALT_INV_RegFile[1][20]~q\ <= NOT \RegFile[1][20]~q\;
\ALT_INV_RegFile[2][20]~q\ <= NOT \RegFile[2][20]~q\;
\ALT_INV_Mux102~0_combout\ <= NOT \Mux102~0_combout\;
\ALT_INV_RegFile[7][20]~q\ <= NOT \RegFile[7][20]~q\;
\ALT_INV_RegFile[6][20]~q\ <= NOT \RegFile[6][20]~q\;
\ALT_INV_RegFile[5][20]~q\ <= NOT \RegFile[5][20]~q\;
\ALT_INV_RegFile[4][20]~q\ <= NOT \RegFile[4][20]~q\;
\ALT_INV_Mux103~13_combout\ <= NOT \Mux103~13_combout\;
\ALT_INV_RegFile[3][19]~q\ <= NOT \RegFile[3][19]~q\;
\ALT_INV_RegFile[1][19]~q\ <= NOT \RegFile[1][19]~q\;
\ALT_INV_RegFile[2][19]~q\ <= NOT \RegFile[2][19]~q\;
\ALT_INV_Mux103~0_combout\ <= NOT \Mux103~0_combout\;
\ALT_INV_RegFile[7][19]~q\ <= NOT \RegFile[7][19]~q\;
\ALT_INV_RegFile[6][19]~q\ <= NOT \RegFile[6][19]~q\;
\ALT_INV_RegFile[5][19]~q\ <= NOT \RegFile[5][19]~q\;
\ALT_INV_RegFile[4][19]~q\ <= NOT \RegFile[4][19]~q\;
\ALT_INV_Mux104~13_combout\ <= NOT \Mux104~13_combout\;
\ALT_INV_RegFile[3][18]~q\ <= NOT \RegFile[3][18]~q\;
\ALT_INV_RegFile[1][18]~q\ <= NOT \RegFile[1][18]~q\;
\ALT_INV_RegFile[2][18]~q\ <= NOT \RegFile[2][18]~q\;
\ALT_INV_Mux104~0_combout\ <= NOT \Mux104~0_combout\;
\ALT_INV_RegFile[7][18]~q\ <= NOT \RegFile[7][18]~q\;
\ALT_INV_RegFile[6][18]~q\ <= NOT \RegFile[6][18]~q\;
\ALT_INV_RegFile[5][18]~q\ <= NOT \RegFile[5][18]~q\;
\ALT_INV_RegFile[4][18]~q\ <= NOT \RegFile[4][18]~q\;
\ALT_INV_Mux105~13_combout\ <= NOT \Mux105~13_combout\;
\ALT_INV_RegFile[3][17]~q\ <= NOT \RegFile[3][17]~q\;
\ALT_INV_RegFile[1][17]~q\ <= NOT \RegFile[1][17]~q\;
\ALT_INV_RegFile[2][17]~q\ <= NOT \RegFile[2][17]~q\;
\ALT_INV_Mux105~0_combout\ <= NOT \Mux105~0_combout\;
\ALT_INV_RegFile[7][17]~q\ <= NOT \RegFile[7][17]~q\;
\ALT_INV_RegFile[6][17]~q\ <= NOT \RegFile[6][17]~q\;
\ALT_INV_RegFile[5][17]~q\ <= NOT \RegFile[5][17]~q\;
\ALT_INV_RegFile[4][17]~q\ <= NOT \RegFile[4][17]~q\;
\ALT_INV_Mux106~13_combout\ <= NOT \Mux106~13_combout\;
\ALT_INV_RegFile[3][16]~q\ <= NOT \RegFile[3][16]~q\;
\ALT_INV_RegFile[1][16]~q\ <= NOT \RegFile[1][16]~q\;
\ALT_INV_RegFile[2][16]~q\ <= NOT \RegFile[2][16]~q\;
\ALT_INV_Mux106~0_combout\ <= NOT \Mux106~0_combout\;
\ALT_INV_RegFile[7][16]~q\ <= NOT \RegFile[7][16]~q\;
\ALT_INV_RegFile[6][16]~q\ <= NOT \RegFile[6][16]~q\;
\ALT_INV_RegFile[5][16]~q\ <= NOT \RegFile[5][16]~q\;
\ALT_INV_RegFile[4][16]~q\ <= NOT \RegFile[4][16]~q\;
\ALT_INV_Mux115~13_combout\ <= NOT \Mux115~13_combout\;
\ALT_INV_RegFile[3][7]~q\ <= NOT \RegFile[3][7]~q\;
\ALT_INV_RegFile[1][7]~q\ <= NOT \RegFile[1][7]~q\;
\ALT_INV_RegFile[2][7]~q\ <= NOT \RegFile[2][7]~q\;
\ALT_INV_Mux115~0_combout\ <= NOT \Mux115~0_combout\;
\ALT_INV_RegFile[7][7]~q\ <= NOT \RegFile[7][7]~q\;
\ALT_INV_RegFile[6][7]~q\ <= NOT \RegFile[6][7]~q\;
\ALT_INV_RegFile[5][7]~q\ <= NOT \RegFile[5][7]~q\;
\ALT_INV_RegFile[4][7]~q\ <= NOT \RegFile[4][7]~q\;
\ALT_INV_Mux107~13_combout\ <= NOT \Mux107~13_combout\;
\ALT_INV_RegFile[3][15]~q\ <= NOT \RegFile[3][15]~q\;
\ALT_INV_RegFile[1][15]~q\ <= NOT \RegFile[1][15]~q\;
\ALT_INV_RegFile[2][15]~q\ <= NOT \RegFile[2][15]~q\;
\ALT_INV_Mux107~0_combout\ <= NOT \Mux107~0_combout\;
\ALT_INV_RegFile[7][15]~q\ <= NOT \RegFile[7][15]~q\;
\ALT_INV_RegFile[6][15]~q\ <= NOT \RegFile[6][15]~q\;
\ALT_INV_RegFile[5][15]~q\ <= NOT \RegFile[5][15]~q\;
\ALT_INV_RegFile[4][15]~q\ <= NOT \RegFile[4][15]~q\;
\ALT_INV_Mux91~13_combout\ <= NOT \Mux91~13_combout\;
\ALT_INV_RegFile[3][31]~q\ <= NOT \RegFile[3][31]~q\;
\ALT_INV_RegFile[1][31]~q\ <= NOT \RegFile[1][31]~q\;
\ALT_INV_RegFile[2][31]~q\ <= NOT \RegFile[2][31]~q\;
\ALT_INV_Mux91~0_combout\ <= NOT \Mux91~0_combout\;
\ALT_INV_RegFile[7][31]~q\ <= NOT \RegFile[7][31]~q\;
\ALT_INV_RegFile[6][31]~q\ <= NOT \RegFile[6][31]~q\;
\ALT_INV_RegFile[5][31]~q\ <= NOT \RegFile[5][31]~q\;
\ALT_INV_RegFile[4][31]~q\ <= NOT \RegFile[4][31]~q\;
\ALT_INV_Mux116~13_combout\ <= NOT \Mux116~13_combout\;
\ALT_INV_RegFile[3][6]~q\ <= NOT \RegFile[3][6]~q\;
\ALT_INV_RegFile[1][6]~q\ <= NOT \RegFile[1][6]~q\;
\ALT_INV_RegFile[2][6]~q\ <= NOT \RegFile[2][6]~q\;
\ALT_INV_Mux116~0_combout\ <= NOT \Mux116~0_combout\;
\ALT_INV_RegFile[7][6]~q\ <= NOT \RegFile[7][6]~q\;
\ALT_INV_RegFile[6][6]~q\ <= NOT \RegFile[6][6]~q\;
\ALT_INV_RegFile[5][6]~q\ <= NOT \RegFile[5][6]~q\;
\ALT_INV_RegFile[4][6]~q\ <= NOT \RegFile[4][6]~q\;
\ALT_INV_Mux108~13_combout\ <= NOT \Mux108~13_combout\;
\ALT_INV_RegFile[3][14]~q\ <= NOT \RegFile[3][14]~q\;
\ALT_INV_RegFile[1][14]~q\ <= NOT \RegFile[1][14]~q\;
\ALT_INV_RegFile[2][14]~q\ <= NOT \RegFile[2][14]~q\;
\ALT_INV_Mux108~0_combout\ <= NOT \Mux108~0_combout\;
\ALT_INV_RegFile[7][14]~q\ <= NOT \RegFile[7][14]~q\;
\ALT_INV_RegFile[6][14]~q\ <= NOT \RegFile[6][14]~q\;
\ALT_INV_RegFile[5][14]~q\ <= NOT \RegFile[5][14]~q\;
\ALT_INV_RegFile[4][14]~q\ <= NOT \RegFile[4][14]~q\;
\ALT_INV_Mux92~13_combout\ <= NOT \Mux92~13_combout\;
\ALT_INV_RegFile[3][30]~q\ <= NOT \RegFile[3][30]~q\;
\ALT_INV_RegFile[1][30]~q\ <= NOT \RegFile[1][30]~q\;
\ALT_INV_RegFile[2][30]~q\ <= NOT \RegFile[2][30]~q\;
\ALT_INV_Mux92~0_combout\ <= NOT \Mux92~0_combout\;
\ALT_INV_RegFile[7][30]~q\ <= NOT \RegFile[7][30]~q\;
\ALT_INV_RegFile[6][30]~q\ <= NOT \RegFile[6][30]~q\;
\ALT_INV_RegFile[5][30]~q\ <= NOT \RegFile[5][30]~q\;
\ALT_INV_RegFile[4][30]~q\ <= NOT \RegFile[4][30]~q\;
\ALT_INV_Mux117~13_combout\ <= NOT \Mux117~13_combout\;
\ALT_INV_RegFile[3][5]~q\ <= NOT \RegFile[3][5]~q\;
\ALT_INV_RegFile[1][5]~q\ <= NOT \RegFile[1][5]~q\;
\ALT_INV_RegFile[2][5]~q\ <= NOT \RegFile[2][5]~q\;
\ALT_INV_Mux117~0_combout\ <= NOT \Mux117~0_combout\;
\ALT_INV_RegFile[7][5]~q\ <= NOT \RegFile[7][5]~q\;
\ALT_INV_RegFile[6][5]~q\ <= NOT \RegFile[6][5]~q\;
\ALT_INV_RegFile[5][5]~q\ <= NOT \RegFile[5][5]~q\;
\ALT_INV_RegFile[4][5]~q\ <= NOT \RegFile[4][5]~q\;
\ALT_INV_Mux109~13_combout\ <= NOT \Mux109~13_combout\;
\ALT_INV_RegFile[3][13]~q\ <= NOT \RegFile[3][13]~q\;
\ALT_INV_RegFile[1][13]~q\ <= NOT \RegFile[1][13]~q\;
\ALT_INV_RegFile[2][13]~q\ <= NOT \RegFile[2][13]~q\;
\ALT_INV_Mux109~0_combout\ <= NOT \Mux109~0_combout\;
\ALT_INV_RegFile[7][13]~q\ <= NOT \RegFile[7][13]~q\;
\ALT_INV_RegFile[6][13]~q\ <= NOT \RegFile[6][13]~q\;
\ALT_INV_RegFile[5][13]~q\ <= NOT \RegFile[5][13]~q\;
\ALT_INV_RegFile[4][13]~q\ <= NOT \RegFile[4][13]~q\;
\ALT_INV_Mux93~13_combout\ <= NOT \Mux93~13_combout\;
\ALT_INV_RegFile[3][29]~q\ <= NOT \RegFile[3][29]~q\;
\ALT_INV_RegFile[1][29]~q\ <= NOT \RegFile[1][29]~q\;
\ALT_INV_RegFile[2][29]~q\ <= NOT \RegFile[2][29]~q\;
\ALT_INV_Mux93~0_combout\ <= NOT \Mux93~0_combout\;
\ALT_INV_RegFile[7][29]~q\ <= NOT \RegFile[7][29]~q\;
\ALT_INV_RegFile[6][29]~q\ <= NOT \RegFile[6][29]~q\;
\ALT_INV_RegFile[5][29]~q\ <= NOT \RegFile[5][29]~q\;
\ALT_INV_RegFile[4][29]~q\ <= NOT \RegFile[4][29]~q\;
\ALT_INV_Mux118~13_combout\ <= NOT \Mux118~13_combout\;
\ALT_INV_RegFile[3][4]~q\ <= NOT \RegFile[3][4]~q\;
\ALT_INV_RegFile[1][4]~q\ <= NOT \RegFile[1][4]~q\;
\ALT_INV_RegFile[2][4]~q\ <= NOT \RegFile[2][4]~q\;
\ALT_INV_Mux118~0_combout\ <= NOT \Mux118~0_combout\;
\ALT_INV_RegFile[7][4]~q\ <= NOT \RegFile[7][4]~q\;
\ALT_INV_RegFile[6][4]~q\ <= NOT \RegFile[6][4]~q\;
\ALT_INV_RegFile[5][4]~q\ <= NOT \RegFile[5][4]~q\;
\ALT_INV_RegFile[4][4]~q\ <= NOT \RegFile[4][4]~q\;
\ALT_INV_Mux110~13_combout\ <= NOT \Mux110~13_combout\;
\ALT_INV_RegFile[3][12]~q\ <= NOT \RegFile[3][12]~q\;
\ALT_INV_RegFile[1][12]~q\ <= NOT \RegFile[1][12]~q\;
\ALT_INV_RegFile[2][12]~q\ <= NOT \RegFile[2][12]~q\;
\ALT_INV_Mux110~0_combout\ <= NOT \Mux110~0_combout\;
\ALT_INV_RegFile[7][12]~q\ <= NOT \RegFile[7][12]~q\;
\ALT_INV_RegFile[6][12]~q\ <= NOT \RegFile[6][12]~q\;
\ALT_INV_RegFile[5][12]~q\ <= NOT \RegFile[5][12]~q\;
\ALT_INV_RegFile[4][12]~q\ <= NOT \RegFile[4][12]~q\;
\ALT_INV_Mux94~13_combout\ <= NOT \Mux94~13_combout\;
\ALT_INV_RegFile[3][28]~q\ <= NOT \RegFile[3][28]~q\;
\ALT_INV_RegFile[1][28]~q\ <= NOT \RegFile[1][28]~q\;
\ALT_INV_RegFile[2][28]~q\ <= NOT \RegFile[2][28]~q\;
\ALT_INV_Mux94~0_combout\ <= NOT \Mux94~0_combout\;
\ALT_INV_RegFile[7][28]~q\ <= NOT \RegFile[7][28]~q\;
\ALT_INV_RegFile[6][28]~q\ <= NOT \RegFile[6][28]~q\;
\ALT_INV_RegFile[5][28]~q\ <= NOT \RegFile[5][28]~q\;
\ALT_INV_RegFile[4][28]~q\ <= NOT \RegFile[4][28]~q\;
\ALT_INV_Mux119~13_combout\ <= NOT \Mux119~13_combout\;
\ALT_INV_RegFile[3][3]~q\ <= NOT \RegFile[3][3]~q\;
\ALT_INV_RegFile[1][3]~q\ <= NOT \RegFile[1][3]~q\;
\ALT_INV_RegFile[2][3]~q\ <= NOT \RegFile[2][3]~q\;
\ALT_INV_Mux119~0_combout\ <= NOT \Mux119~0_combout\;
\ALT_INV_RegFile[7][3]~q\ <= NOT \RegFile[7][3]~q\;
\ALT_INV_RegFile[6][3]~q\ <= NOT \RegFile[6][3]~q\;
\ALT_INV_RegFile[5][3]~q\ <= NOT \RegFile[5][3]~q\;
\ALT_INV_RegFile[4][3]~q\ <= NOT \RegFile[4][3]~q\;
\ALT_INV_Mux111~13_combout\ <= NOT \Mux111~13_combout\;
\ALT_INV_RegFile[3][11]~q\ <= NOT \RegFile[3][11]~q\;
\ALT_INV_RegFile[1][11]~q\ <= NOT \RegFile[1][11]~q\;
\ALT_INV_RegFile[2][11]~q\ <= NOT \RegFile[2][11]~q\;
\ALT_INV_Mux111~0_combout\ <= NOT \Mux111~0_combout\;
\ALT_INV_RegFile[7][11]~q\ <= NOT \RegFile[7][11]~q\;
\ALT_INV_RegFile[6][11]~q\ <= NOT \RegFile[6][11]~q\;
\ALT_INV_RegFile[5][11]~q\ <= NOT \RegFile[5][11]~q\;
\ALT_INV_RegFile[4][11]~q\ <= NOT \RegFile[4][11]~q\;
\ALT_INV_Mux95~13_combout\ <= NOT \Mux95~13_combout\;
\ALT_INV_RegFile[3][27]~q\ <= NOT \RegFile[3][27]~q\;
\ALT_INV_RegFile[1][27]~q\ <= NOT \RegFile[1][27]~q\;
\ALT_INV_RegFile[2][27]~q\ <= NOT \RegFile[2][27]~q\;
\ALT_INV_Mux95~0_combout\ <= NOT \Mux95~0_combout\;
\ALT_INV_RegFile[7][27]~q\ <= NOT \RegFile[7][27]~q\;
\ALT_INV_RegFile[6][27]~q\ <= NOT \RegFile[6][27]~q\;
\ALT_INV_RegFile[5][27]~q\ <= NOT \RegFile[5][27]~q\;
\ALT_INV_RegFile[4][27]~q\ <= NOT \RegFile[4][27]~q\;
\ALT_INV_Mux120~13_combout\ <= NOT \Mux120~13_combout\;
\ALT_INV_RegFile[3][2]~q\ <= NOT \RegFile[3][2]~q\;
\ALT_INV_RegFile[1][2]~q\ <= NOT \RegFile[1][2]~q\;
\ALT_INV_RegFile[2][2]~q\ <= NOT \RegFile[2][2]~q\;
\ALT_INV_Mux120~0_combout\ <= NOT \Mux120~0_combout\;
\ALT_INV_RegFile[7][2]~q\ <= NOT \RegFile[7][2]~q\;
\ALT_INV_RegFile[6][2]~q\ <= NOT \RegFile[6][2]~q\;
\ALT_INV_RegFile[5][2]~q\ <= NOT \RegFile[5][2]~q\;
\ALT_INV_RegFile[4][2]~q\ <= NOT \RegFile[4][2]~q\;
\ALT_INV_Mux112~13_combout\ <= NOT \Mux112~13_combout\;
\ALT_INV_RegFile[3][10]~q\ <= NOT \RegFile[3][10]~q\;
\ALT_INV_RegFile[1][10]~q\ <= NOT \RegFile[1][10]~q\;
\ALT_INV_RegFile[2][10]~q\ <= NOT \RegFile[2][10]~q\;
\ALT_INV_Mux112~0_combout\ <= NOT \Mux112~0_combout\;
\ALT_INV_RegFile[7][10]~q\ <= NOT \RegFile[7][10]~q\;
\ALT_INV_RegFile[6][10]~q\ <= NOT \RegFile[6][10]~q\;
\ALT_INV_RegFile[5][10]~q\ <= NOT \RegFile[5][10]~q\;
\ALT_INV_RegFile[4][10]~q\ <= NOT \RegFile[4][10]~q\;
\ALT_INV_Mux96~13_combout\ <= NOT \Mux96~13_combout\;
\ALT_INV_RegFile[3][26]~q\ <= NOT \RegFile[3][26]~q\;
\ALT_INV_RegFile[1][26]~q\ <= NOT \RegFile[1][26]~q\;
\ALT_INV_RegFile[2][26]~q\ <= NOT \RegFile[2][26]~q\;
\ALT_INV_Mux96~0_combout\ <= NOT \Mux96~0_combout\;
\ALT_INV_RegFile[7][26]~q\ <= NOT \RegFile[7][26]~q\;
\ALT_INV_RegFile[6][26]~q\ <= NOT \RegFile[6][26]~q\;
\ALT_INV_RegFile[5][26]~q\ <= NOT \RegFile[5][26]~q\;
\ALT_INV_RegFile[4][26]~q\ <= NOT \RegFile[4][26]~q\;
\ALT_INV_Mux121~13_combout\ <= NOT \Mux121~13_combout\;
\ALT_INV_RegFile[3][1]~q\ <= NOT \RegFile[3][1]~q\;
\ALT_INV_RegFile[1][1]~q\ <= NOT \RegFile[1][1]~q\;
\ALT_INV_RegFile[2][1]~q\ <= NOT \RegFile[2][1]~q\;
\ALT_INV_Mux121~0_combout\ <= NOT \Mux121~0_combout\;
\ALT_INV_RegFile[7][1]~q\ <= NOT \RegFile[7][1]~q\;
\ALT_INV_RegFile[6][1]~q\ <= NOT \RegFile[6][1]~q\;
\ALT_INV_RegFile[5][1]~q\ <= NOT \RegFile[5][1]~q\;
\ALT_INV_RegFile[4][1]~q\ <= NOT \RegFile[4][1]~q\;
\ALT_INV_Mux113~13_combout\ <= NOT \Mux113~13_combout\;
\ALT_INV_RegFile[3][9]~q\ <= NOT \RegFile[3][9]~q\;
\ALT_INV_RegFile[1][9]~q\ <= NOT \RegFile[1][9]~q\;
\ALT_INV_RegFile[2][9]~q\ <= NOT \RegFile[2][9]~q\;
\ALT_INV_Mux113~0_combout\ <= NOT \Mux113~0_combout\;
\ALT_INV_RegFile[7][9]~q\ <= NOT \RegFile[7][9]~q\;
\ALT_INV_RegFile[6][9]~q\ <= NOT \RegFile[6][9]~q\;
\ALT_INV_RegFile[5][9]~q\ <= NOT \RegFile[5][9]~q\;
\ALT_INV_RegFile[4][9]~q\ <= NOT \RegFile[4][9]~q\;
\ALT_INV_Mux97~13_combout\ <= NOT \Mux97~13_combout\;
\ALT_INV_RegFile[3][25]~q\ <= NOT \RegFile[3][25]~q\;
\ALT_INV_RegFile[1][25]~q\ <= NOT \RegFile[1][25]~q\;
\ALT_INV_RegFile[2][25]~q\ <= NOT \RegFile[2][25]~q\;
\ALT_INV_Mux97~0_combout\ <= NOT \Mux97~0_combout\;
\ALT_INV_RegFile[7][25]~q\ <= NOT \RegFile[7][25]~q\;
\ALT_INV_RegFile[6][25]~q\ <= NOT \RegFile[6][25]~q\;
\ALT_INV_RegFile[5][25]~q\ <= NOT \RegFile[5][25]~q\;
\ALT_INV_RegFile[4][25]~q\ <= NOT \RegFile[4][25]~q\;
\ALT_INV_Mux122~13_combout\ <= NOT \Mux122~13_combout\;
\ALT_INV_RegFile[3][0]~q\ <= NOT \RegFile[3][0]~q\;
\ALT_INV_RegFile[1][0]~q\ <= NOT \RegFile[1][0]~q\;
\ALT_INV_RegFile[2][0]~q\ <= NOT \RegFile[2][0]~q\;
\ALT_INV_Mux122~0_combout\ <= NOT \Mux122~0_combout\;
\ALT_INV_RegFile[7][0]~q\ <= NOT \RegFile[7][0]~q\;
\ALT_INV_RegFile[6][0]~q\ <= NOT \RegFile[6][0]~q\;
\ALT_INV_RegFile[5][0]~q\ <= NOT \RegFile[5][0]~q\;
\ALT_INV_RegFile[4][0]~q\ <= NOT \RegFile[4][0]~q\;
\ALT_INV_Mux114~13_combout\ <= NOT \Mux114~13_combout\;
\ALT_INV_RegFile[3][8]~q\ <= NOT \RegFile[3][8]~q\;
\ALT_INV_RegFile[1][8]~q\ <= NOT \RegFile[1][8]~q\;
\ALT_INV_RegFile[2][8]~q\ <= NOT \RegFile[2][8]~q\;
\ALT_INV_Mux114~0_combout\ <= NOT \Mux114~0_combout\;
\ALT_INV_RegFile[7][8]~q\ <= NOT \RegFile[7][8]~q\;
\ALT_INV_RegFile[6][8]~q\ <= NOT \RegFile[6][8]~q\;
\ALT_INV_RegFile[5][8]~q\ <= NOT \RegFile[5][8]~q\;
\ALT_INV_RegFile[4][8]~q\ <= NOT \RegFile[4][8]~q\;
\ALT_INV_Mux98~13_combout\ <= NOT \Mux98~13_combout\;
\ALT_INV_R.curInst\(24) <= NOT \R.curInst\(24);
\ALT_INV_R.curInst\(23) <= NOT \R.curInst\(23);
\ALT_INV_RegFile[3][24]~q\ <= NOT \RegFile[3][24]~q\;
\ALT_INV_RegFile[1][24]~q\ <= NOT \RegFile[1][24]~q\;
\ALT_INV_RegFile[2][24]~q\ <= NOT \RegFile[2][24]~q\;
\ALT_INV_Mux98~0_combout\ <= NOT \Mux98~0_combout\;
\ALT_INV_R.curInst\(21) <= NOT \R.curInst\(21);
\ALT_INV_R.curInst\(20) <= NOT \R.curInst\(20);
\ALT_INV_RegFile[7][24]~q\ <= NOT \RegFile[7][24]~q\;
\ALT_INV_RegFile[6][24]~q\ <= NOT \RegFile[6][24]~q\;
\ALT_INV_RegFile[5][24]~q\ <= NOT \RegFile[5][24]~q\;
\ALT_INV_RegFile[4][24]~q\ <= NOT \RegFile[4][24]~q\;
\ALT_INV_R.curInst\(22) <= NOT \R.curInst\(22);
\ALT_INV_Mux162~0_combout\ <= NOT \Mux162~0_combout\;
\ALT_INV_Mux221~0_combout\ <= NOT \Mux221~0_combout\;
\ALT_INV_Mux222~0_combout\ <= NOT \Mux222~0_combout\;
\ALT_INV_R.curInst\(12) <= NOT \R.curInst\(12);
\ALT_INV_R.curInst\(14) <= NOT \R.curInst\(14);
\ALT_INV_R.curInst\(13) <= NOT \R.curInst\(13);
\ALT_INV_R.aluRes\(31) <= NOT \R.aluRes\(31);
\ALT_INV_Selector1~2_combout\ <= NOT \Selector1~2_combout\;
\ALT_INV_Selector1~1_combout\ <= NOT \Selector1~1_combout\;
\ALT_INV_ShiftLeft0~56_combout\ <= NOT \ShiftLeft0~56_combout\;
\ALT_INV_R.aluRes\(30) <= NOT \R.aluRes\(30);
\ALT_INV_Selector2~2_combout\ <= NOT \Selector2~2_combout\;
\ALT_INV_Selector2~1_combout\ <= NOT \Selector2~1_combout\;
\ALT_INV_Selector2~0_combout\ <= NOT \Selector2~0_combout\;
\ALT_INV_ShiftLeft0~54_combout\ <= NOT \ShiftLeft0~54_combout\;
\ALT_INV_R.aluRes\(29) <= NOT \R.aluRes\(29);
\ALT_INV_Selector3~2_combout\ <= NOT \Selector3~2_combout\;
\ALT_INV_Selector3~1_combout\ <= NOT \Selector3~1_combout\;
\ALT_INV_Selector3~0_combout\ <= NOT \Selector3~0_combout\;
\ALT_INV_ShiftLeft0~52_combout\ <= NOT \ShiftLeft0~52_combout\;
\ALT_INV_R.aluRes\(28) <= NOT \R.aluRes\(28);
\ALT_INV_Selector4~1_combout\ <= NOT \Selector4~1_combout\;
\ALT_INV_Selector4~0_combout\ <= NOT \Selector4~0_combout\;
\ALT_INV_ShiftLeft0~50_combout\ <= NOT \ShiftLeft0~50_combout\;
\ALT_INV_Selector20~5_combout\ <= NOT \Selector20~5_combout\;
\ALT_INV_R.aluRes\(27) <= NOT \R.aluRes\(27);
\ALT_INV_Selector5~4_combout\ <= NOT \Selector5~4_combout\;
\ALT_INV_Selector5~3_combout\ <= NOT \Selector5~3_combout\;
\ALT_INV_Selector5~2_combout\ <= NOT \Selector5~2_combout\;
\ALT_INV_Selector5~1_combout\ <= NOT \Selector5~1_combout\;
\ALT_INV_ShiftLeft0~48_combout\ <= NOT \ShiftLeft0~48_combout\;
\ALT_INV_Selector5~0_combout\ <= NOT \Selector5~0_combout\;
\ALT_INV_R.aluRes\(26) <= NOT \R.aluRes\(26);
\ALT_INV_Selector6~2_combout\ <= NOT \Selector6~2_combout\;
\ALT_INV_Selector6~1_combout\ <= NOT \Selector6~1_combout\;
\ALT_INV_Selector6~0_combout\ <= NOT \Selector6~0_combout\;
\ALT_INV_ShiftLeft0~46_combout\ <= NOT \ShiftLeft0~46_combout\;
\ALT_INV_ShiftLeft0~44_combout\ <= NOT \ShiftLeft0~44_combout\;
\ALT_INV_R.aluRes\(25) <= NOT \R.aluRes\(25);
\ALT_INV_Selector7~3_combout\ <= NOT \Selector7~3_combout\;
\ALT_INV_Selector7~2_combout\ <= NOT \Selector7~2_combout\;
\ALT_INV_Selector7~1_combout\ <= NOT \Selector7~1_combout\;
\ALT_INV_ShiftLeft0~43_combout\ <= NOT \ShiftLeft0~43_combout\;
\ALT_INV_Selector7~0_combout\ <= NOT \Selector7~0_combout\;
\ALT_INV_ShiftRight1~55_combout\ <= NOT \ShiftRight1~55_combout\;
\ALT_INV_R.aluRes\(24) <= NOT \R.aluRes\(24);
\ALT_INV_Selector8~4_combout\ <= NOT \Selector8~4_combout\;
\ALT_INV_Selector8~3_combout\ <= NOT \Selector8~3_combout\;
\ALT_INV_Selector8~2_combout\ <= NOT \Selector8~2_combout\;
\ALT_INV_Selector8~1_combout\ <= NOT \Selector8~1_combout\;
\ALT_INV_Selector8~0_combout\ <= NOT \Selector8~0_combout\;
\ALT_INV_ShiftLeft0~41_combout\ <= NOT \ShiftLeft0~41_combout\;
\ALT_INV_R.aluRes\(23) <= NOT \R.aluRes\(23);
\ALT_INV_Selector9~5_combout\ <= NOT \Selector9~5_combout\;
\ALT_INV_Selector9~4_combout\ <= NOT \Selector9~4_combout\;
\ALT_INV_Selector9~3_combout\ <= NOT \Selector9~3_combout\;
\ALT_INV_Selector9~2_combout\ <= NOT \Selector9~2_combout\;
\ALT_INV_Selector9~1_combout\ <= NOT \Selector9~1_combout\;
\ALT_INV_ShiftLeft0~39_combout\ <= NOT \ShiftLeft0~39_combout\;
\ALT_INV_Selector9~0_combout\ <= NOT \Selector9~0_combout\;
\ALT_INV_ShiftRight0~12_combout\ <= NOT \ShiftRight0~12_combout\;
\ALT_INV_R.aluRes\(22) <= NOT \R.aluRes\(22);
\ALT_INV_Selector10~4_combout\ <= NOT \Selector10~4_combout\;
\ALT_INV_Selector10~3_combout\ <= NOT \Selector10~3_combout\;
\ALT_INV_Selector10~2_combout\ <= NOT \Selector10~2_combout\;
\ALT_INV_Selector10~1_combout\ <= NOT \Selector10~1_combout\;
\ALT_INV_ShiftLeft0~37_combout\ <= NOT \ShiftLeft0~37_combout\;
\ALT_INV_Selector10~0_combout\ <= NOT \Selector10~0_combout\;
\ALT_INV_R.aluRes\(21) <= NOT \R.aluRes\(21);
\ALT_INV_Selector11~5_combout\ <= NOT \Selector11~5_combout\;
\ALT_INV_Selector11~4_combout\ <= NOT \Selector11~4_combout\;
\ALT_INV_Selector11~3_combout\ <= NOT \Selector11~3_combout\;
\ALT_INV_Selector11~2_combout\ <= NOT \Selector11~2_combout\;
\ALT_INV_Selector11~1_combout\ <= NOT \Selector11~1_combout\;
\ALT_INV_ShiftLeft0~35_combout\ <= NOT \ShiftLeft0~35_combout\;
\ALT_INV_Selector11~0_combout\ <= NOT \Selector11~0_combout\;
\ALT_INV_vAluRes~17_combout\ <= NOT \vAluRes~17_combout\;
\ALT_INV_R.aluRes\(20) <= NOT \R.aluRes\(20);
\ALT_INV_Selector12~5_combout\ <= NOT \Selector12~5_combout\;
\ALT_INV_Selector12~4_combout\ <= NOT \Selector12~4_combout\;
\ALT_INV_Selector12~3_combout\ <= NOT \Selector12~3_combout\;
\ALT_INV_Selector12~1_combout\ <= NOT \Selector12~1_combout\;
\ALT_INV_ShiftLeft0~33_combout\ <= NOT \ShiftLeft0~33_combout\;
\ALT_INV_Selector12~0_combout\ <= NOT \Selector12~0_combout\;
\ALT_INV_R.aluRes\(19) <= NOT \R.aluRes\(19);
\ALT_INV_Selector13~1_combout\ <= NOT \Selector13~1_combout\;
\ALT_INV_Selector13~0_combout\ <= NOT \Selector13~0_combout\;
\ALT_INV_ShiftLeft0~31_combout\ <= NOT \ShiftLeft0~31_combout\;
\ALT_INV_R.aluRes\(18) <= NOT \R.aluRes\(18);
\ALT_INV_Selector14~3_combout\ <= NOT \Selector14~3_combout\;
\ALT_INV_Selector14~2_combout\ <= NOT \Selector14~2_combout\;
\ALT_INV_Selector14~1_combout\ <= NOT \Selector14~1_combout\;
\ALT_INV_Selector14~0_combout\ <= NOT \Selector14~0_combout\;
\ALT_INV_ShiftLeft0~29_combout\ <= NOT \ShiftLeft0~29_combout\;
\ALT_INV_R.aluRes\(17) <= NOT \R.aluRes\(17);
\ALT_INV_Selector15~4_combout\ <= NOT \Selector15~4_combout\;
\ALT_INV_Selector15~3_combout\ <= NOT \Selector15~3_combout\;
\ALT_INV_ShiftLeft0~27_combout\ <= NOT \ShiftLeft0~27_combout\;
\ALT_INV_Selector15~1_combout\ <= NOT \Selector15~1_combout\;
\ALT_INV_Selector15~0_combout\ <= NOT \Selector15~0_combout\;
\ALT_INV_R.aluRes\(16) <= NOT \R.aluRes\(16);
\ALT_INV_Selector16~4_combout\ <= NOT \Selector16~4_combout\;
\ALT_INV_Selector16~3_combout\ <= NOT \Selector16~3_combout\;
\ALT_INV_Selector16~2_combout\ <= NOT \Selector16~2_combout\;
\ALT_INV_ShiftLeft0~25_combout\ <= NOT \ShiftLeft0~25_combout\;
\ALT_INV_R.aluRes\(15) <= NOT \R.aluRes\(15);
\ALT_INV_Selector17~3_combout\ <= NOT \Selector17~3_combout\;
\ALT_INV_Selector17~2_combout\ <= NOT \Selector17~2_combout\;
\ALT_INV_Selector17~1_combout\ <= NOT \Selector17~1_combout\;
\ALT_INV_ShiftRight1~54_combout\ <= NOT \ShiftRight1~54_combout\;
\ALT_INV_ShiftLeft0~23_combout\ <= NOT \ShiftLeft0~23_combout\;
\ALT_INV_R.aluRes\(14) <= NOT \R.aluRes\(14);
\ALT_INV_Selector18~4_combout\ <= NOT \Selector18~4_combout\;
\ALT_INV_Selector18~3_combout\ <= NOT \Selector18~3_combout\;
\ALT_INV_Selector18~2_combout\ <= NOT \Selector18~2_combout\;
\ALT_INV_Selector18~0_combout\ <= NOT \Selector18~0_combout\;
\ALT_INV_ShiftRight1~53_combout\ <= NOT \ShiftRight1~53_combout\;
\ALT_INV_ShiftLeft0~21_combout\ <= NOT \ShiftLeft0~21_combout\;
\ALT_INV_R.aluRes\(13) <= NOT \R.aluRes\(13);
\ALT_INV_Selector19~3_combout\ <= NOT \Selector19~3_combout\;
\ALT_INV_Selector19~2_combout\ <= NOT \Selector19~2_combout\;
\ALT_INV_Selector19~1_combout\ <= NOT \Selector19~1_combout\;
\ALT_INV_ShiftRight1~52_combout\ <= NOT \ShiftRight1~52_combout\;
\ALT_INV_ShiftLeft0~19_combout\ <= NOT \ShiftLeft0~19_combout\;
\ALT_INV_R.aluRes\(12) <= NOT \R.aluRes\(12);
\ALT_INV_Selector20~4_combout\ <= NOT \Selector20~4_combout\;
\ALT_INV_Selector20~3_combout\ <= NOT \Selector20~3_combout\;
\ALT_INV_Selector20~2_combout\ <= NOT \Selector20~2_combout\;
\ALT_INV_ShiftRight1~51_combout\ <= NOT \ShiftRight1~51_combout\;
\ALT_INV_Selector20~1_combout\ <= NOT \Selector20~1_combout\;
\ALT_INV_ShiftLeft0~17_combout\ <= NOT \ShiftLeft0~17_combout\;
\ALT_INV_R.aluRes\(11) <= NOT \R.aluRes\(11);
\ALT_INV_Selector21~3_combout\ <= NOT \Selector21~3_combout\;
\ALT_INV_Selector21~2_combout\ <= NOT \Selector21~2_combout\;
\ALT_INV_Selector21~1_combout\ <= NOT \Selector21~1_combout\;
\ALT_INV_ShiftRight1~50_combout\ <= NOT \ShiftRight1~50_combout\;
\ALT_INV_Selector21~0_combout\ <= NOT \Selector21~0_combout\;
\ALT_INV_ShiftLeft0~15_combout\ <= NOT \ShiftLeft0~15_combout\;
\ALT_INV_vAluRes~10_combout\ <= NOT \vAluRes~10_combout\;
\ALT_INV_R.aluRes\(10) <= NOT \R.aluRes\(10);
\ALT_INV_Selector22~4_combout\ <= NOT \Selector22~4_combout\;
\ALT_INV_ShiftRight1~49_combout\ <= NOT \ShiftRight1~49_combout\;
\ALT_INV_Selector22~3_combout\ <= NOT \Selector22~3_combout\;
\ALT_INV_Selector22~2_combout\ <= NOT \Selector22~2_combout\;
\ALT_INV_R.aluRes\(9) <= NOT \R.aluRes\(9);
\ALT_INV_Selector23~5_combout\ <= NOT \Selector23~5_combout\;
\ALT_INV_Selector23~4_combout\ <= NOT \Selector23~4_combout\;
\ALT_INV_ShiftRight1~47_combout\ <= NOT \ShiftRight1~47_combout\;
\ALT_INV_Selector23~2_combout\ <= NOT \Selector23~2_combout\;
\ALT_INV_Selector23~1_combout\ <= NOT \Selector23~1_combout\;
\ALT_INV_Selector23~0_combout\ <= NOT \Selector23~0_combout\;
\ALT_INV_vAluRes~8_combout\ <= NOT \vAluRes~8_combout\;
\ALT_INV_R.aluRes\(8) <= NOT \R.aluRes\(8);
\ALT_INV_Selector24~3_combout\ <= NOT \Selector24~3_combout\;
\ALT_INV_ShiftRight1~46_combout\ <= NOT \ShiftRight1~46_combout\;
\ALT_INV_ShiftRight0~10_combout\ <= NOT \ShiftRight0~10_combout\;
\ALT_INV_ShiftLeft0~11_combout\ <= NOT \ShiftLeft0~11_combout\;
\ALT_INV_Selector24~1_combout\ <= NOT \Selector24~1_combout\;
\ALT_INV_vAluRes~7_combout\ <= NOT \vAluRes~7_combout\;
\ALT_INV_R.aluRes\(7) <= NOT \R.aluRes\(7);
\ALT_INV_Selector25~4_combout\ <= NOT \Selector25~4_combout\;
\ALT_INV_ShiftRight1~45_combout\ <= NOT \ShiftRight1~45_combout\;
\ALT_INV_Selector25~2_combout\ <= NOT \Selector25~2_combout\;
\ALT_INV_Selector25~1_combout\ <= NOT \Selector25~1_combout\;
\ALT_INV_vAluRes~6_combout\ <= NOT \vAluRes~6_combout\;
\ALT_INV_R.aluRes\(6) <= NOT \R.aluRes\(6);
\ALT_INV_Selector26~3_combout\ <= NOT \Selector26~3_combout\;
\ALT_INV_ShiftRight1~44_combout\ <= NOT \ShiftRight1~44_combout\;
\ALT_INV_ShiftRight0~9_combout\ <= NOT \ShiftRight0~9_combout\;
\ALT_INV_Selector26~1_combout\ <= NOT \Selector26~1_combout\;
\ALT_INV_Selector26~0_combout\ <= NOT \Selector26~0_combout\;
\ALT_INV_ShiftRight1~43_combout\ <= NOT \ShiftRight1~43_combout\;
\ALT_INV_vAluRes~5_combout\ <= NOT \vAluRes~5_combout\;
\ALT_INV_R.aluRes\(5) <= NOT \R.aluRes\(5);
\ALT_INV_Selector27~4_combout\ <= NOT \Selector27~4_combout\;
\ALT_INV_Selector27~3_combout\ <= NOT \Selector27~3_combout\;
\ALT_INV_ShiftRight1~42_combout\ <= NOT \ShiftRight1~42_combout\;
\ALT_INV_ShiftRight0~8_combout\ <= NOT \ShiftRight0~8_combout\;
\ALT_INV_Selector27~1_combout\ <= NOT \Selector27~1_combout\;
\ALT_INV_ShiftRight1~41_combout\ <= NOT \ShiftRight1~41_combout\;
\ALT_INV_vAluRes~4_combout\ <= NOT \vAluRes~4_combout\;
\ALT_INV_R.aluRes\(4) <= NOT \R.aluRes\(4);
\ALT_INV_Selector28~3_combout\ <= NOT \Selector28~3_combout\;
\ALT_INV_Selector28~2_combout\ <= NOT \Selector28~2_combout\;
\ALT_INV_ShiftRight1~40_combout\ <= NOT \ShiftRight1~40_combout\;
\ALT_INV_ShiftRight0~6_combout\ <= NOT \ShiftRight0~6_combout\;
\ALT_INV_Selector28~0_combout\ <= NOT \Selector28~0_combout\;
\ALT_INV_ShiftRight1~39_combout\ <= NOT \ShiftRight1~39_combout\;
\ALT_INV_vAluRes~3_combout\ <= NOT \vAluRes~3_combout\;
\ALT_INV_R.aluRes\(3) <= NOT \R.aluRes\(3);
\ALT_INV_Selector29~3_combout\ <= NOT \Selector29~3_combout\;
\ALT_INV_Selector29~2_combout\ <= NOT \Selector29~2_combout\;
\ALT_INV_Selector29~1_combout\ <= NOT \Selector29~1_combout\;
\ALT_INV_ShiftRight1~38_combout\ <= NOT \ShiftRight1~38_combout\;
\ALT_INV_ShiftRight1~33_combout\ <= NOT \ShiftRight1~33_combout\;
\ALT_INV_ShiftRight0~5_combout\ <= NOT \ShiftRight0~5_combout\;
\ALT_INV_vAluRes~2_combout\ <= NOT \vAluRes~2_combout\;
\ALT_INV_R.aluRes\(2) <= NOT \R.aluRes\(2);
\ALT_INV_Selector30~3_combout\ <= NOT \Selector30~3_combout\;
\ALT_INV_Selector30~2_combout\ <= NOT \Selector30~2_combout\;
\ALT_INV_ShiftRight0~3_combout\ <= NOT \ShiftRight0~3_combout\;
\ALT_INV_Selector30~0_combout\ <= NOT \Selector30~0_combout\;
\ALT_INV_ShiftRight1~29_combout\ <= NOT \ShiftRight1~29_combout\;
\ALT_INV_ShiftRight1~24_combout\ <= NOT \ShiftRight1~24_combout\;
\ALT_INV_ShiftRight1~20_combout\ <= NOT \ShiftRight1~20_combout\;
\ALT_INV_vAluRes~1_combout\ <= NOT \vAluRes~1_combout\;
\ALT_INV_R.aluRes\(1) <= NOT \R.aluRes\(1);
\ALT_INV_Selector31~4_combout\ <= NOT \Selector31~4_combout\;
\ALT_INV_Selector31~3_combout\ <= NOT \Selector31~3_combout\;
\ALT_INV_Selector31~1_combout\ <= NOT \Selector31~1_combout\;
\ALT_INV_ShiftRight1~19_combout\ <= NOT \ShiftRight1~19_combout\;
\ALT_INV_ShiftRight0~1_combout\ <= NOT \ShiftRight0~1_combout\;
\ALT_INV_ShiftRight1~14_combout\ <= NOT \ShiftRight1~14_combout\;
\ALT_INV_vAluRes~0_combout\ <= NOT \vAluRes~0_combout\;
\ALT_INV_R.aluRes\(0) <= NOT \R.aluRes\(0);
\ALT_INV_Selector32~7_combout\ <= NOT \Selector32~7_combout\;
\ALT_INV_R.aluOp.ALUOpAnd~q\ <= NOT \R.aluOp.ALUOpAnd~q\;
\ALT_INV_R.aluOp.ALUOpOr~q\ <= NOT \R.aluOp.ALUOpOr~q\;
\ALT_INV_R.aluOp.ALUOpSLL~q\ <= NOT \R.aluOp.ALUOpSLL~q\;
\ALT_INV_R.aluOp.ALUOpSub~q\ <= NOT \R.aluOp.ALUOpSub~q\;
\ALT_INV_Selector32~2_combout\ <= NOT \Selector32~2_combout\;
\ALT_INV_R.aluOp.ALUOpAdd~q\ <= NOT \R.aluOp.ALUOpAdd~q\;
\ALT_INV_R.aluOp.ALUOpXor~q\ <= NOT \R.aluOp.ALUOpXor~q\;
\ALT_INV_ShiftRight1~9_combout\ <= NOT \ShiftRight1~9_combout\;
\ALT_INV_ShiftRight1~4_combout\ <= NOT \ShiftRight1~4_combout\;
\ALT_INV_R.aluOp.ALUOpSRA~q\ <= NOT \R.aluOp.ALUOpSRA~q\;
\ALT_INV_R.aluOp.ALUOpSRL~q\ <= NOT \R.aluOp.ALUOpSRL~q\;
\ALT_INV_Selector32~1_combout\ <= NOT \Selector32~1_combout\;
\ALT_INV_LessThan1~38_combout\ <= NOT \LessThan1~38_combout\;
\ALT_INV_LessThan1~37_combout\ <= NOT \LessThan1~37_combout\;
\ALT_INV_R.aluData2\(29) <= NOT \R.aluData2\(29);
\ALT_INV_R.aluData1\(29) <= NOT \R.aluData1\(29);
\ALT_INV_R.aluData2\(30) <= NOT \R.aluData2\(30);
\ALT_INV_R.aluData1\(30) <= NOT \R.aluData1\(30);
\ALT_INV_R.aluData2\(31) <= NOT \R.aluData2\(31);
\ALT_INV_R.aluData1\(31) <= NOT \R.aluData1\(31);
\ALT_INV_LessThan1~36_combout\ <= NOT \LessThan1~36_combout\;
\ALT_INV_LessThan1~35_combout\ <= NOT \LessThan1~35_combout\;
\ALT_INV_LessThan1~33_combout\ <= NOT \LessThan1~33_combout\;
\ALT_INV_LessThan1~32_combout\ <= NOT \LessThan1~32_combout\;
\ALT_INV_LessThan1~31_combout\ <= NOT \LessThan1~31_combout\;
\ALT_INV_R.aluData2\(22) <= NOT \R.aluData2\(22);
\ALT_INV_R.aluData1\(22) <= NOT \R.aluData1\(22);
\ALT_INV_R.aluData2\(23) <= NOT \R.aluData2\(23);
\ALT_INV_R.aluData1\(23) <= NOT \R.aluData1\(23);
\ALT_INV_R.aluData2\(24) <= NOT \R.aluData2\(24);
\ALT_INV_R.aluData1\(24) <= NOT \R.aluData1\(24);
\ALT_INV_R.aluData2\(26) <= NOT \R.aluData2\(26);
\ALT_INV_R.aluData1\(26) <= NOT \R.aluData1\(26);
\ALT_INV_R.aluData2\(27) <= NOT \R.aluData2\(27);
\ALT_INV_R.aluData1\(27) <= NOT \R.aluData1\(27);
\ALT_INV_R.aluData2\(28) <= NOT \R.aluData2\(28);
\ALT_INV_R.aluData1\(28) <= NOT \R.aluData1\(28);
\ALT_INV_R.aluData2\(25) <= NOT \R.aluData2\(25);
\ALT_INV_R.aluData1\(25) <= NOT \R.aluData1\(25);
\ALT_INV_LessThan1~27_combout\ <= NOT \LessThan1~27_combout\;
\ALT_INV_LessThan1~26_combout\ <= NOT \LessThan1~26_combout\;
\ALT_INV_LessThan1~23_combout\ <= NOT \LessThan1~23_combout\;
\ALT_INV_LessThan1~19_combout\ <= NOT \LessThan1~19_combout\;
\ALT_INV_LessThan1~17_combout\ <= NOT \LessThan1~17_combout\;
\ALT_INV_LessThan1~13_combout\ <= NOT \LessThan1~13_combout\;
\ALT_INV_R.aluData1\(4) <= NOT \R.aluData1\(4);
\ALT_INV_R.aluData1\(5) <= NOT \R.aluData1\(5);
\ALT_INV_R.aluData2\(4) <= NOT \R.aluData2\(4);
\ALT_INV_R.aluData1\(2) <= NOT \R.aluData1\(2);
\ALT_INV_R.aluData1\(3) <= NOT \R.aluData1\(3);
\ALT_INV_R.aluData2\(2) <= NOT \R.aluData2\(2);
\ALT_INV_R.aluData2\(3) <= NOT \R.aluData2\(3);
\ALT_INV_R.aluData2\(1) <= NOT \R.aluData2\(1);
\ALT_INV_R.aluData2\(0) <= NOT \R.aluData2\(0);
\ALT_INV_LessThan1~6_combout\ <= NOT \LessThan1~6_combout\;
\ALT_INV_R.aluData2\(12) <= NOT \R.aluData2\(12);
\ALT_INV_R.aluData1\(12) <= NOT \R.aluData1\(12);
\ALT_INV_R.aluData2\(13) <= NOT \R.aluData2\(13);
\ALT_INV_R.aluData1\(13) <= NOT \R.aluData1\(13);
\ALT_INV_R.aluData2\(11) <= NOT \R.aluData2\(11);
\ALT_INV_R.aluData1\(11) <= NOT \R.aluData1\(11);
\ALT_INV_R.aluData2\(15) <= NOT \R.aluData2\(15);
\ALT_INV_R.aluData1\(15) <= NOT \R.aluData1\(15);
\ALT_INV_R.aluData2\(18) <= NOT \R.aluData2\(18);
\ALT_INV_R.aluData1\(18) <= NOT \R.aluData1\(18);
\ALT_INV_R.aluData2\(19) <= NOT \R.aluData2\(19);
\ALT_INV_R.aluData1\(19) <= NOT \R.aluData1\(19);
\ALT_INV_R.aluData2\(20) <= NOT \R.aluData2\(20);
\ALT_INV_R.aluData1\(20) <= NOT \R.aluData1\(20);
\ALT_INV_R.aluData2\(21) <= NOT \R.aluData2\(21);
\ALT_INV_R.aluData1\(21) <= NOT \R.aluData1\(21);
\ALT_INV_Selector32~0_combout\ <= NOT \Selector32~0_combout\;
\ALT_INV_R.aluOp.ALUOpSLT~q\ <= NOT \R.aluOp.ALUOpSLT~q\;
\ALT_INV_R.aluOp.ALUOpSLTU~q\ <= NOT \R.aluOp.ALUOpSLTU~q\;
\ALT_INV_Comb~0_combout\ <= NOT \Comb~0_combout\;
\ALT_INV_R.ctrlState.WriteReg~q\ <= NOT \R.ctrlState.WriteReg~q\;
\ALT_INV_R.ctrlState.Wait1~q\ <= NOT \R.ctrlState.Wait1~q\;
\ALT_INV_R.curPC\(1) <= NOT \R.curPC\(1);
\ALT_INV_vAluRes~60_combout\ <= NOT \vAluRes~60_combout\;
\ALT_INV_vAluRes~56_combout\ <= NOT \vAluRes~56_combout\;
\ALT_INV_vAluRes~52_combout\ <= NOT \vAluRes~52_combout\;
\ALT_INV_Selector7~5_combout\ <= NOT \Selector7~5_combout\;
\ALT_INV_Mux98~26_combout\ <= NOT \Mux98~26_combout\;
\ALT_INV_Mux114~26_combout\ <= NOT \Mux114~26_combout\;
\ALT_INV_Mux122~26_combout\ <= NOT \Mux122~26_combout\;
\ALT_INV_Mux97~26_combout\ <= NOT \Mux97~26_combout\;
\ALT_INV_Mux113~26_combout\ <= NOT \Mux113~26_combout\;
\ALT_INV_Mux121~26_combout\ <= NOT \Mux121~26_combout\;
\ALT_INV_Mux96~26_combout\ <= NOT \Mux96~26_combout\;
\ALT_INV_Mux112~26_combout\ <= NOT \Mux112~26_combout\;
\ALT_INV_Mux120~26_combout\ <= NOT \Mux120~26_combout\;
\ALT_INV_Mux95~26_combout\ <= NOT \Mux95~26_combout\;
\ALT_INV_Mux111~26_combout\ <= NOT \Mux111~26_combout\;
\ALT_INV_Mux119~26_combout\ <= NOT \Mux119~26_combout\;
\ALT_INV_Mux94~26_combout\ <= NOT \Mux94~26_combout\;
\ALT_INV_Mux110~26_combout\ <= NOT \Mux110~26_combout\;
\ALT_INV_Mux118~26_combout\ <= NOT \Mux118~26_combout\;
\ALT_INV_Mux93~26_combout\ <= NOT \Mux93~26_combout\;
\ALT_INV_Mux109~26_combout\ <= NOT \Mux109~26_combout\;
\ALT_INV_Mux117~26_combout\ <= NOT \Mux117~26_combout\;
\ALT_INV_Mux92~26_combout\ <= NOT \Mux92~26_combout\;
\ALT_INV_Mux108~26_combout\ <= NOT \Mux108~26_combout\;
\ALT_INV_Mux116~26_combout\ <= NOT \Mux116~26_combout\;
\ALT_INV_Mux91~26_combout\ <= NOT \Mux91~26_combout\;
\ALT_INV_Mux107~26_combout\ <= NOT \Mux107~26_combout\;
\ALT_INV_Mux115~26_combout\ <= NOT \Mux115~26_combout\;
\ALT_INV_Mux106~26_combout\ <= NOT \Mux106~26_combout\;
\ALT_INV_Mux105~26_combout\ <= NOT \Mux105~26_combout\;
\ALT_INV_Mux104~26_combout\ <= NOT \Mux104~26_combout\;
\ALT_INV_Mux103~26_combout\ <= NOT \Mux103~26_combout\;
\ALT_INV_Mux102~26_combout\ <= NOT \Mux102~26_combout\;
\ALT_INV_Mux101~26_combout\ <= NOT \Mux101~26_combout\;
\ALT_INV_Mux100~26_combout\ <= NOT \Mux100~26_combout\;
\ALT_INV_Mux99~26_combout\ <= NOT \Mux99~26_combout\;
\ALT_INV_Mux19~0_combout\ <= NOT \Mux19~0_combout\;
\ALT_INV_Mux69~26_combout\ <= NOT \Mux69~26_combout\;
\ALT_INV_Mux70~26_combout\ <= NOT \Mux70~26_combout\;
\ALT_INV_Mux71~26_combout\ <= NOT \Mux71~26_combout\;
\ALT_INV_Mux72~26_combout\ <= NOT \Mux72~26_combout\;
\ALT_INV_Mux73~26_combout\ <= NOT \Mux73~26_combout\;
\ALT_INV_Mux74~26_combout\ <= NOT \Mux74~26_combout\;
\ALT_INV_Mux75~26_combout\ <= NOT \Mux75~26_combout\;
\ALT_INV_Mux76~26_combout\ <= NOT \Mux76~26_combout\;
\ALT_INV_Mux79~26_combout\ <= NOT \Mux79~26_combout\;
\ALT_INV_Mux80~26_combout\ <= NOT \Mux80~26_combout\;
\ALT_INV_Mux77~26_combout\ <= NOT \Mux77~26_combout\;
\ALT_INV_Mux78~26_combout\ <= NOT \Mux78~26_combout\;
\ALT_INV_Mux81~26_combout\ <= NOT \Mux81~26_combout\;
\ALT_INV_Mux82~26_combout\ <= NOT \Mux82~26_combout\;
\ALT_INV_Mux83~26_combout\ <= NOT \Mux83~26_combout\;
\ALT_INV_Mux84~26_combout\ <= NOT \Mux84~26_combout\;
\ALT_INV_Mux90~26_combout\ <= NOT \Mux90~26_combout\;
\ALT_INV_Mux89~26_combout\ <= NOT \Mux89~26_combout\;
\ALT_INV_Mux87~26_combout\ <= NOT \Mux87~26_combout\;
\ALT_INV_Mux88~26_combout\ <= NOT \Mux88~26_combout\;
\ALT_INV_Mux85~26_combout\ <= NOT \Mux85~26_combout\;
\ALT_INV_Mux86~26_combout\ <= NOT \Mux86~26_combout\;
\ALT_INV_Mux65~26_combout\ <= NOT \Mux65~26_combout\;
\ALT_INV_Mux62~26_combout\ <= NOT \Mux62~26_combout\;
\ALT_INV_Mux63~26_combout\ <= NOT \Mux63~26_combout\;
\ALT_INV_Mux64~26_combout\ <= NOT \Mux64~26_combout\;
\ALT_INV_Mux66~26_combout\ <= NOT \Mux66~26_combout\;
\ALT_INV_Mux67~26_combout\ <= NOT \Mux67~26_combout\;
\ALT_INV_Mux68~26_combout\ <= NOT \Mux68~26_combout\;
\ALT_INV_Mux59~26_combout\ <= NOT \Mux59~26_combout\;
\ALT_INV_Mux60~26_combout\ <= NOT \Mux60~26_combout\;
\ALT_INV_Mux61~26_combout\ <= NOT \Mux61~26_combout\;
\ALT_INV_Add1~129_sumout\ <= NOT \Add1~129_sumout\;
\ALT_INV_Add2~129_sumout\ <= NOT \Add2~129_sumout\;
\ALT_INV_R.csrRead~q\ <= NOT \R.csrRead~q\;
\ALT_INV_R.memToReg~q\ <= NOT \R.memToReg~q\;
\ALT_INV_Mux61~22_combout\ <= NOT \Mux61~22_combout\;
\ALT_INV_Mux61~18_combout\ <= NOT \Mux61~18_combout\;
\ALT_INV_Mux61~14_combout\ <= NOT \Mux61~14_combout\;
\ALT_INV_Mux60~22_combout\ <= NOT \Mux60~22_combout\;
\ALT_INV_Mux60~18_combout\ <= NOT \Mux60~18_combout\;
\ALT_INV_Mux60~14_combout\ <= NOT \Mux60~14_combout\;
\ALT_INV_Mux59~22_combout\ <= NOT \Mux59~22_combout\;
\ALT_INV_Mux59~18_combout\ <= NOT \Mux59~18_combout\;
\ALT_INV_Mux59~14_combout\ <= NOT \Mux59~14_combout\;
\ALT_INV_Mux68~22_combout\ <= NOT \Mux68~22_combout\;
\ALT_INV_Mux68~18_combout\ <= NOT \Mux68~18_combout\;
\ALT_INV_Mux68~14_combout\ <= NOT \Mux68~14_combout\;
\ALT_INV_Mux67~22_combout\ <= NOT \Mux67~22_combout\;
\ALT_INV_Mux67~18_combout\ <= NOT \Mux67~18_combout\;
\ALT_INV_Mux67~14_combout\ <= NOT \Mux67~14_combout\;
\ALT_INV_Mux66~22_combout\ <= NOT \Mux66~22_combout\;
\ALT_INV_Mux66~18_combout\ <= NOT \Mux66~18_combout\;
\ALT_INV_Mux66~14_combout\ <= NOT \Mux66~14_combout\;
\ALT_INV_Mux64~22_combout\ <= NOT \Mux64~22_combout\;
\ALT_INV_Mux64~18_combout\ <= NOT \Mux64~18_combout\;
\ALT_INV_Mux64~14_combout\ <= NOT \Mux64~14_combout\;
\ALT_INV_Mux63~22_combout\ <= NOT \Mux63~22_combout\;
\ALT_INV_Mux63~18_combout\ <= NOT \Mux63~18_combout\;
\ALT_INV_Mux63~14_combout\ <= NOT \Mux63~14_combout\;
\ALT_INV_Mux62~22_combout\ <= NOT \Mux62~22_combout\;
\ALT_INV_Mux62~18_combout\ <= NOT \Mux62~18_combout\;
\ALT_INV_Mux62~14_combout\ <= NOT \Mux62~14_combout\;
\ALT_INV_Mux65~22_combout\ <= NOT \Mux65~22_combout\;
\ALT_INV_Mux65~18_combout\ <= NOT \Mux65~18_combout\;
\ALT_INV_Mux65~14_combout\ <= NOT \Mux65~14_combout\;
\ALT_INV_Mux86~22_combout\ <= NOT \Mux86~22_combout\;
\ALT_INV_Mux86~18_combout\ <= NOT \Mux86~18_combout\;
\ALT_INV_Mux86~14_combout\ <= NOT \Mux86~14_combout\;
\ALT_INV_Mux85~22_combout\ <= NOT \Mux85~22_combout\;
\ALT_INV_Mux85~18_combout\ <= NOT \Mux85~18_combout\;
\ALT_INV_Mux85~14_combout\ <= NOT \Mux85~14_combout\;
\ALT_INV_Mux88~22_combout\ <= NOT \Mux88~22_combout\;
\ALT_INV_Mux88~18_combout\ <= NOT \Mux88~18_combout\;
\ALT_INV_Mux88~14_combout\ <= NOT \Mux88~14_combout\;
\ALT_INV_Mux87~22_combout\ <= NOT \Mux87~22_combout\;
\ALT_INV_Mux87~18_combout\ <= NOT \Mux87~18_combout\;
\ALT_INV_Mux87~14_combout\ <= NOT \Mux87~14_combout\;
\ALT_INV_Mux89~22_combout\ <= NOT \Mux89~22_combout\;
\ALT_INV_Mux89~18_combout\ <= NOT \Mux89~18_combout\;
\ALT_INV_Mux89~14_combout\ <= NOT \Mux89~14_combout\;
\ALT_INV_Mux90~22_combout\ <= NOT \Mux90~22_combout\;
\ALT_INV_Mux90~18_combout\ <= NOT \Mux90~18_combout\;
\ALT_INV_Mux90~14_combout\ <= NOT \Mux90~14_combout\;
\ALT_INV_Mux84~22_combout\ <= NOT \Mux84~22_combout\;
\ALT_INV_Mux84~18_combout\ <= NOT \Mux84~18_combout\;
\ALT_INV_Mux84~14_combout\ <= NOT \Mux84~14_combout\;
\ALT_INV_Mux83~22_combout\ <= NOT \Mux83~22_combout\;
\ALT_INV_Mux83~18_combout\ <= NOT \Mux83~18_combout\;
\ALT_INV_Mux83~14_combout\ <= NOT \Mux83~14_combout\;
\ALT_INV_Mux82~22_combout\ <= NOT \Mux82~22_combout\;
\ALT_INV_Mux82~18_combout\ <= NOT \Mux82~18_combout\;
\ALT_INV_Mux82~14_combout\ <= NOT \Mux82~14_combout\;
\ALT_INV_Mux81~22_combout\ <= NOT \Mux81~22_combout\;
\ALT_INV_Mux81~18_combout\ <= NOT \Mux81~18_combout\;
\ALT_INV_Mux81~14_combout\ <= NOT \Mux81~14_combout\;
\ALT_INV_Mux78~22_combout\ <= NOT \Mux78~22_combout\;
\ALT_INV_Mux78~18_combout\ <= NOT \Mux78~18_combout\;
\ALT_INV_Mux78~14_combout\ <= NOT \Mux78~14_combout\;
\ALT_INV_Mux77~22_combout\ <= NOT \Mux77~22_combout\;
\ALT_INV_Mux77~18_combout\ <= NOT \Mux77~18_combout\;
\ALT_INV_Mux77~14_combout\ <= NOT \Mux77~14_combout\;
\ALT_INV_Mux80~22_combout\ <= NOT \Mux80~22_combout\;
\ALT_INV_Mux80~18_combout\ <= NOT \Mux80~18_combout\;
\ALT_INV_Mux80~14_combout\ <= NOT \Mux80~14_combout\;
\ALT_INV_Mux79~22_combout\ <= NOT \Mux79~22_combout\;
\ALT_INV_Mux79~18_combout\ <= NOT \Mux79~18_combout\;
\ALT_INV_Mux79~14_combout\ <= NOT \Mux79~14_combout\;
\ALT_INV_Mux76~22_combout\ <= NOT \Mux76~22_combout\;
\ALT_INV_Mux76~18_combout\ <= NOT \Mux76~18_combout\;
\ALT_INV_Mux76~14_combout\ <= NOT \Mux76~14_combout\;
\ALT_INV_Mux75~22_combout\ <= NOT \Mux75~22_combout\;
\ALT_INV_Mux75~18_combout\ <= NOT \Mux75~18_combout\;
\ALT_INV_Mux75~14_combout\ <= NOT \Mux75~14_combout\;
\ALT_INV_Mux74~22_combout\ <= NOT \Mux74~22_combout\;
\ALT_INV_Mux74~18_combout\ <= NOT \Mux74~18_combout\;
\ALT_INV_Mux74~14_combout\ <= NOT \Mux74~14_combout\;
\ALT_INV_Mux73~22_combout\ <= NOT \Mux73~22_combout\;
\ALT_INV_Mux73~18_combout\ <= NOT \Mux73~18_combout\;
\ALT_INV_Mux73~14_combout\ <= NOT \Mux73~14_combout\;
\ALT_INV_Mux72~22_combout\ <= NOT \Mux72~22_combout\;
\ALT_INV_Mux72~18_combout\ <= NOT \Mux72~18_combout\;
\ALT_INV_Mux72~14_combout\ <= NOT \Mux72~14_combout\;
\ALT_INV_Mux71~22_combout\ <= NOT \Mux71~22_combout\;
\ALT_INV_Mux71~18_combout\ <= NOT \Mux71~18_combout\;
\ALT_INV_Mux71~14_combout\ <= NOT \Mux71~14_combout\;
\ALT_INV_Mux70~22_combout\ <= NOT \Mux70~22_combout\;
\ALT_INV_Mux70~18_combout\ <= NOT \Mux70~18_combout\;
\ALT_INV_Mux70~14_combout\ <= NOT \Mux70~14_combout\;
\ALT_INV_Mux69~22_combout\ <= NOT \Mux69~22_combout\;
\ALT_INV_Mux69~18_combout\ <= NOT \Mux69~18_combout\;
\ALT_INV_Mux69~14_combout\ <= NOT \Mux69~14_combout\;
\ALT_INV_Mux99~22_combout\ <= NOT \Mux99~22_combout\;
\ALT_INV_Mux99~18_combout\ <= NOT \Mux99~18_combout\;
\ALT_INV_Mux99~14_combout\ <= NOT \Mux99~14_combout\;
\ALT_INV_R.regWriteData\(23) <= NOT \R.regWriteData\(23);
\ALT_INV_Mux100~22_combout\ <= NOT \Mux100~22_combout\;
\ALT_INV_Mux100~18_combout\ <= NOT \Mux100~18_combout\;
\ALT_INV_Mux100~14_combout\ <= NOT \Mux100~14_combout\;
\ALT_INV_R.regWriteData\(22) <= NOT \R.regWriteData\(22);
\ALT_INV_Mux101~22_combout\ <= NOT \Mux101~22_combout\;
\ALT_INV_Mux101~18_combout\ <= NOT \Mux101~18_combout\;
\ALT_INV_Mux101~14_combout\ <= NOT \Mux101~14_combout\;
\ALT_INV_R.regWriteData\(21) <= NOT \R.regWriteData\(21);
\ALT_INV_Mux102~22_combout\ <= NOT \Mux102~22_combout\;
\ALT_INV_Mux102~18_combout\ <= NOT \Mux102~18_combout\;
\ALT_INV_Mux102~14_combout\ <= NOT \Mux102~14_combout\;
\ALT_INV_R.regWriteData\(20) <= NOT \R.regWriteData\(20);
\ALT_INV_Mux103~22_combout\ <= NOT \Mux103~22_combout\;
\ALT_INV_Mux103~18_combout\ <= NOT \Mux103~18_combout\;
\ALT_INV_Mux103~14_combout\ <= NOT \Mux103~14_combout\;
\ALT_INV_R.regWriteData\(19) <= NOT \R.regWriteData\(19);
\ALT_INV_Mux104~22_combout\ <= NOT \Mux104~22_combout\;
\ALT_INV_Mux104~18_combout\ <= NOT \Mux104~18_combout\;
\ALT_INV_Mux104~14_combout\ <= NOT \Mux104~14_combout\;
\ALT_INV_R.regWriteData\(18) <= NOT \R.regWriteData\(18);
\ALT_INV_Mux105~22_combout\ <= NOT \Mux105~22_combout\;
\ALT_INV_Mux105~18_combout\ <= NOT \Mux105~18_combout\;
\ALT_INV_Mux105~14_combout\ <= NOT \Mux105~14_combout\;
\ALT_INV_R.regWriteData\(17) <= NOT \R.regWriteData\(17);
\ALT_INV_Mux106~22_combout\ <= NOT \Mux106~22_combout\;
\ALT_INV_Mux106~18_combout\ <= NOT \Mux106~18_combout\;
\ALT_INV_Mux106~14_combout\ <= NOT \Mux106~14_combout\;
\ALT_INV_R.regWriteData\(16) <= NOT \R.regWriteData\(16);
\ALT_INV_Mux115~22_combout\ <= NOT \Mux115~22_combout\;
\ALT_INV_Mux115~18_combout\ <= NOT \Mux115~18_combout\;
\ALT_INV_Mux115~14_combout\ <= NOT \Mux115~14_combout\;
\ALT_INV_R.regWriteData\(7) <= NOT \R.regWriteData\(7);
\ALT_INV_Mux107~22_combout\ <= NOT \Mux107~22_combout\;
\ALT_INV_Mux107~18_combout\ <= NOT \Mux107~18_combout\;
\ALT_INV_Mux107~14_combout\ <= NOT \Mux107~14_combout\;
\ALT_INV_R.regWriteData\(15) <= NOT \R.regWriteData\(15);
\ALT_INV_Mux91~22_combout\ <= NOT \Mux91~22_combout\;
\ALT_INV_Mux91~18_combout\ <= NOT \Mux91~18_combout\;
\ALT_INV_Mux91~14_combout\ <= NOT \Mux91~14_combout\;
\ALT_INV_R.regWriteData\(31) <= NOT \R.regWriteData\(31);
\ALT_INV_Mux116~22_combout\ <= NOT \Mux116~22_combout\;
\ALT_INV_Mux116~18_combout\ <= NOT \Mux116~18_combout\;
\ALT_INV_Mux116~14_combout\ <= NOT \Mux116~14_combout\;
\ALT_INV_R.regWriteData\(6) <= NOT \R.regWriteData\(6);
\ALT_INV_Mux108~22_combout\ <= NOT \Mux108~22_combout\;
\ALT_INV_Mux108~18_combout\ <= NOT \Mux108~18_combout\;
\ALT_INV_Mux108~14_combout\ <= NOT \Mux108~14_combout\;
\ALT_INV_R.regWriteData\(14) <= NOT \R.regWriteData\(14);
\ALT_INV_Mux92~22_combout\ <= NOT \Mux92~22_combout\;
\ALT_INV_Mux92~18_combout\ <= NOT \Mux92~18_combout\;
\ALT_INV_Mux92~14_combout\ <= NOT \Mux92~14_combout\;
\ALT_INV_R.regWriteData\(30) <= NOT \R.regWriteData\(30);
\ALT_INV_Mux117~22_combout\ <= NOT \Mux117~22_combout\;
\ALT_INV_Mux117~18_combout\ <= NOT \Mux117~18_combout\;
\ALT_INV_Mux117~14_combout\ <= NOT \Mux117~14_combout\;
\ALT_INV_R.regWriteData\(5) <= NOT \R.regWriteData\(5);
\ALT_INV_Mux109~22_combout\ <= NOT \Mux109~22_combout\;
\ALT_INV_Mux109~18_combout\ <= NOT \Mux109~18_combout\;
\ALT_INV_Mux109~14_combout\ <= NOT \Mux109~14_combout\;
\ALT_INV_R.regWriteData\(13) <= NOT \R.regWriteData\(13);
\ALT_INV_Mux93~22_combout\ <= NOT \Mux93~22_combout\;
\ALT_INV_Mux93~18_combout\ <= NOT \Mux93~18_combout\;
\ALT_INV_Mux93~14_combout\ <= NOT \Mux93~14_combout\;
\ALT_INV_R.regWriteData\(29) <= NOT \R.regWriteData\(29);
\ALT_INV_Mux118~22_combout\ <= NOT \Mux118~22_combout\;
\ALT_INV_Mux118~18_combout\ <= NOT \Mux118~18_combout\;
\ALT_INV_Mux118~14_combout\ <= NOT \Mux118~14_combout\;
\ALT_INV_R.regWriteData\(4) <= NOT \R.regWriteData\(4);
\ALT_INV_Mux110~22_combout\ <= NOT \Mux110~22_combout\;
\ALT_INV_Mux110~18_combout\ <= NOT \Mux110~18_combout\;
\ALT_INV_Mux110~14_combout\ <= NOT \Mux110~14_combout\;
\ALT_INV_R.regWriteData\(12) <= NOT \R.regWriteData\(12);
\ALT_INV_Mux94~22_combout\ <= NOT \Mux94~22_combout\;
\ALT_INV_Mux94~18_combout\ <= NOT \Mux94~18_combout\;
\ALT_INV_Mux94~14_combout\ <= NOT \Mux94~14_combout\;
\ALT_INV_R.regWriteData\(28) <= NOT \R.regWriteData\(28);
\ALT_INV_Mux119~22_combout\ <= NOT \Mux119~22_combout\;
\ALT_INV_Mux119~18_combout\ <= NOT \Mux119~18_combout\;
\ALT_INV_Mux119~14_combout\ <= NOT \Mux119~14_combout\;
\ALT_INV_R.regWriteData\(3) <= NOT \R.regWriteData\(3);
\ALT_INV_Mux111~22_combout\ <= NOT \Mux111~22_combout\;
\ALT_INV_Mux111~18_combout\ <= NOT \Mux111~18_combout\;
\ALT_INV_Mux111~14_combout\ <= NOT \Mux111~14_combout\;
\ALT_INV_R.regWriteData\(11) <= NOT \R.regWriteData\(11);
\ALT_INV_Mux95~22_combout\ <= NOT \Mux95~22_combout\;
\ALT_INV_Mux95~18_combout\ <= NOT \Mux95~18_combout\;
\ALT_INV_Mux95~14_combout\ <= NOT \Mux95~14_combout\;
\ALT_INV_R.regWriteData\(27) <= NOT \R.regWriteData\(27);
\ALT_INV_Mux120~22_combout\ <= NOT \Mux120~22_combout\;
\ALT_INV_Mux120~18_combout\ <= NOT \Mux120~18_combout\;
\ALT_INV_Mux120~14_combout\ <= NOT \Mux120~14_combout\;
\ALT_INV_R.regWriteData\(2) <= NOT \R.regWriteData\(2);
\ALT_INV_Mux112~22_combout\ <= NOT \Mux112~22_combout\;
\ALT_INV_Mux112~18_combout\ <= NOT \Mux112~18_combout\;
\ALT_INV_Mux112~14_combout\ <= NOT \Mux112~14_combout\;
\ALT_INV_R.regWriteData\(10) <= NOT \R.regWriteData\(10);
\ALT_INV_Mux96~22_combout\ <= NOT \Mux96~22_combout\;
\ALT_INV_Mux96~18_combout\ <= NOT \Mux96~18_combout\;
\ALT_INV_Mux96~14_combout\ <= NOT \Mux96~14_combout\;
\ALT_INV_R.regWriteData\(26) <= NOT \R.regWriteData\(26);
\ALT_INV_Mux121~22_combout\ <= NOT \Mux121~22_combout\;
\ALT_INV_Mux121~18_combout\ <= NOT \Mux121~18_combout\;
\ALT_INV_Mux121~14_combout\ <= NOT \Mux121~14_combout\;
\ALT_INV_R.regWriteData\(1) <= NOT \R.regWriteData\(1);
\ALT_INV_Mux113~22_combout\ <= NOT \Mux113~22_combout\;
\ALT_INV_Mux113~18_combout\ <= NOT \Mux113~18_combout\;
\ALT_INV_Mux113~14_combout\ <= NOT \Mux113~14_combout\;
\ALT_INV_R.regWriteData\(9) <= NOT \R.regWriteData\(9);
\ALT_INV_Mux97~22_combout\ <= NOT \Mux97~22_combout\;
\ALT_INV_Mux97~18_combout\ <= NOT \Mux97~18_combout\;
\ALT_INV_Mux97~14_combout\ <= NOT \Mux97~14_combout\;
\ALT_INV_R.regWriteData\(25) <= NOT \R.regWriteData\(25);
\ALT_INV_Mux122~22_combout\ <= NOT \Mux122~22_combout\;
\ALT_INV_Mux122~18_combout\ <= NOT \Mux122~18_combout\;
\ALT_INV_Mux122~14_combout\ <= NOT \Mux122~14_combout\;
\ALT_INV_R.regWriteData\(0) <= NOT \R.regWriteData\(0);
\ALT_INV_Mux114~22_combout\ <= NOT \Mux114~22_combout\;
\ALT_INV_Mux114~18_combout\ <= NOT \Mux114~18_combout\;
\ALT_INV_Mux114~14_combout\ <= NOT \Mux114~14_combout\;
\ALT_INV_R.regWriteData\(8) <= NOT \R.regWriteData\(8);
\ALT_INV_Mux98~22_combout\ <= NOT \Mux98~22_combout\;
\ALT_INV_Mux98~18_combout\ <= NOT \Mux98~18_combout\;
\ALT_INV_Mux98~14_combout\ <= NOT \Mux98~14_combout\;
\ALT_INV_R.regWriteData\(24) <= NOT \R.regWriteData\(24);
\ALT_INV_Mux61~9_combout\ <= NOT \Mux61~9_combout\;
\ALT_INV_Mux61~5_combout\ <= NOT \Mux61~5_combout\;
\ALT_INV_Mux61~1_combout\ <= NOT \Mux61~1_combout\;
\ALT_INV_Mux60~9_combout\ <= NOT \Mux60~9_combout\;
\ALT_INV_Mux60~5_combout\ <= NOT \Mux60~5_combout\;
\ALT_INV_Mux60~1_combout\ <= NOT \Mux60~1_combout\;
\ALT_INV_Mux59~9_combout\ <= NOT \Mux59~9_combout\;
\ALT_INV_Mux59~5_combout\ <= NOT \Mux59~5_combout\;
\ALT_INV_Mux59~1_combout\ <= NOT \Mux59~1_combout\;
\ALT_INV_Mux68~9_combout\ <= NOT \Mux68~9_combout\;
\ALT_INV_Mux68~5_combout\ <= NOT \Mux68~5_combout\;
\ALT_INV_Mux68~1_combout\ <= NOT \Mux68~1_combout\;
\ALT_INV_Mux67~9_combout\ <= NOT \Mux67~9_combout\;
\ALT_INV_Mux67~5_combout\ <= NOT \Mux67~5_combout\;
\ALT_INV_Mux67~1_combout\ <= NOT \Mux67~1_combout\;
\ALT_INV_Mux66~9_combout\ <= NOT \Mux66~9_combout\;
\ALT_INV_Mux66~5_combout\ <= NOT \Mux66~5_combout\;
\ALT_INV_Mux66~1_combout\ <= NOT \Mux66~1_combout\;
\ALT_INV_Mux64~9_combout\ <= NOT \Mux64~9_combout\;
\ALT_INV_Mux64~5_combout\ <= NOT \Mux64~5_combout\;
\ALT_INV_Mux64~1_combout\ <= NOT \Mux64~1_combout\;
\ALT_INV_Mux63~9_combout\ <= NOT \Mux63~9_combout\;
\ALT_INV_Mux63~5_combout\ <= NOT \Mux63~5_combout\;
\ALT_INV_Mux63~1_combout\ <= NOT \Mux63~1_combout\;
\ALT_INV_Mux62~9_combout\ <= NOT \Mux62~9_combout\;
\ALT_INV_Mux62~5_combout\ <= NOT \Mux62~5_combout\;
\ALT_INV_Mux62~1_combout\ <= NOT \Mux62~1_combout\;
\ALT_INV_Mux65~9_combout\ <= NOT \Mux65~9_combout\;
\ALT_INV_Mux65~5_combout\ <= NOT \Mux65~5_combout\;
\ALT_INV_Mux65~1_combout\ <= NOT \Mux65~1_combout\;
\ALT_INV_Mux86~9_combout\ <= NOT \Mux86~9_combout\;
\ALT_INV_Mux86~5_combout\ <= NOT \Mux86~5_combout\;
\ALT_INV_Mux86~1_combout\ <= NOT \Mux86~1_combout\;
\ALT_INV_Mux85~9_combout\ <= NOT \Mux85~9_combout\;
\ALT_INV_Mux85~5_combout\ <= NOT \Mux85~5_combout\;
\ALT_INV_Mux85~1_combout\ <= NOT \Mux85~1_combout\;
\ALT_INV_Mux88~9_combout\ <= NOT \Mux88~9_combout\;
\ALT_INV_Mux88~5_combout\ <= NOT \Mux88~5_combout\;
\ALT_INV_Mux88~1_combout\ <= NOT \Mux88~1_combout\;
\ALT_INV_Mux87~9_combout\ <= NOT \Mux87~9_combout\;
\ALT_INV_Mux87~5_combout\ <= NOT \Mux87~5_combout\;
\ALT_INV_Mux87~1_combout\ <= NOT \Mux87~1_combout\;
\ALT_INV_Mux89~9_combout\ <= NOT \Mux89~9_combout\;
\ALT_INV_Mux89~5_combout\ <= NOT \Mux89~5_combout\;
\ALT_INV_Mux89~1_combout\ <= NOT \Mux89~1_combout\;
\ALT_INV_Mux90~9_combout\ <= NOT \Mux90~9_combout\;
\ALT_INV_Mux90~5_combout\ <= NOT \Mux90~5_combout\;
\ALT_INV_Mux90~1_combout\ <= NOT \Mux90~1_combout\;
\ALT_INV_Mux84~9_combout\ <= NOT \Mux84~9_combout\;
\ALT_INV_Mux84~5_combout\ <= NOT \Mux84~5_combout\;
\ALT_INV_Mux84~1_combout\ <= NOT \Mux84~1_combout\;
\ALT_INV_Mux83~9_combout\ <= NOT \Mux83~9_combout\;
\ALT_INV_Mux83~5_combout\ <= NOT \Mux83~5_combout\;
\ALT_INV_Mux83~1_combout\ <= NOT \Mux83~1_combout\;
\ALT_INV_Mux82~9_combout\ <= NOT \Mux82~9_combout\;
\ALT_INV_Mux82~5_combout\ <= NOT \Mux82~5_combout\;
\ALT_INV_Mux82~1_combout\ <= NOT \Mux82~1_combout\;
\ALT_INV_Mux81~9_combout\ <= NOT \Mux81~9_combout\;
\ALT_INV_Mux81~5_combout\ <= NOT \Mux81~5_combout\;
\ALT_INV_Mux81~1_combout\ <= NOT \Mux81~1_combout\;
\ALT_INV_Mux78~9_combout\ <= NOT \Mux78~9_combout\;
\ALT_INV_Mux78~5_combout\ <= NOT \Mux78~5_combout\;
\ALT_INV_Mux78~1_combout\ <= NOT \Mux78~1_combout\;
\ALT_INV_Mux77~9_combout\ <= NOT \Mux77~9_combout\;
\ALT_INV_Mux77~5_combout\ <= NOT \Mux77~5_combout\;
\ALT_INV_Mux77~1_combout\ <= NOT \Mux77~1_combout\;
\ALT_INV_Mux80~9_combout\ <= NOT \Mux80~9_combout\;
\ALT_INV_Mux80~5_combout\ <= NOT \Mux80~5_combout\;
\ALT_INV_Mux80~1_combout\ <= NOT \Mux80~1_combout\;
\ALT_INV_Mux79~9_combout\ <= NOT \Mux79~9_combout\;
\ALT_INV_Mux79~5_combout\ <= NOT \Mux79~5_combout\;
\ALT_INV_Mux79~1_combout\ <= NOT \Mux79~1_combout\;
\ALT_INV_Mux76~9_combout\ <= NOT \Mux76~9_combout\;
\ALT_INV_Mux76~5_combout\ <= NOT \Mux76~5_combout\;
\ALT_INV_Mux76~1_combout\ <= NOT \Mux76~1_combout\;
\ALT_INV_Mux75~9_combout\ <= NOT \Mux75~9_combout\;
\ALT_INV_Mux75~5_combout\ <= NOT \Mux75~5_combout\;
\ALT_INV_Mux75~1_combout\ <= NOT \Mux75~1_combout\;
\ALT_INV_Mux74~9_combout\ <= NOT \Mux74~9_combout\;
\ALT_INV_Mux74~5_combout\ <= NOT \Mux74~5_combout\;
\ALT_INV_Mux74~1_combout\ <= NOT \Mux74~1_combout\;
\ALT_INV_Mux73~9_combout\ <= NOT \Mux73~9_combout\;
\ALT_INV_Mux73~5_combout\ <= NOT \Mux73~5_combout\;
\ALT_INV_Mux73~1_combout\ <= NOT \Mux73~1_combout\;
\ALT_INV_Mux72~9_combout\ <= NOT \Mux72~9_combout\;
\ALT_INV_Mux72~5_combout\ <= NOT \Mux72~5_combout\;
\ALT_INV_Mux72~1_combout\ <= NOT \Mux72~1_combout\;
\ALT_INV_Mux71~9_combout\ <= NOT \Mux71~9_combout\;
\ALT_INV_Mux71~5_combout\ <= NOT \Mux71~5_combout\;
\ALT_INV_Mux71~1_combout\ <= NOT \Mux71~1_combout\;
\ALT_INV_Mux70~9_combout\ <= NOT \Mux70~9_combout\;
\ALT_INV_Mux70~5_combout\ <= NOT \Mux70~5_combout\;
\ALT_INV_Mux70~1_combout\ <= NOT \Mux70~1_combout\;
\ALT_INV_Mux69~9_combout\ <= NOT \Mux69~9_combout\;
\ALT_INV_Mux69~5_combout\ <= NOT \Mux69~5_combout\;
\ALT_INV_Mux69~1_combout\ <= NOT \Mux69~1_combout\;
\ALT_INV_Add3~125_sumout\ <= NOT \Add3~125_sumout\;
\ALT_INV_Add3~121_sumout\ <= NOT \Add3~121_sumout\;
\ALT_INV_Add3~117_sumout\ <= NOT \Add3~117_sumout\;
\ALT_INV_Add3~113_sumout\ <= NOT \Add3~113_sumout\;
\ALT_INV_Add3~109_sumout\ <= NOT \Add3~109_sumout\;
\ALT_INV_Add3~105_sumout\ <= NOT \Add3~105_sumout\;
\ALT_INV_Add3~101_sumout\ <= NOT \Add3~101_sumout\;
\ALT_INV_Add3~97_sumout\ <= NOT \Add3~97_sumout\;
\ALT_INV_Add3~93_sumout\ <= NOT \Add3~93_sumout\;
\ALT_INV_Add3~89_sumout\ <= NOT \Add3~89_sumout\;
\ALT_INV_Add0~77_sumout\ <= NOT \Add0~77_sumout\;
\ALT_INV_Add3~85_sumout\ <= NOT \Add3~85_sumout\;
\ALT_INV_Add0~73_sumout\ <= NOT \Add0~73_sumout\;
\ALT_INV_Add3~81_sumout\ <= NOT \Add3~81_sumout\;
\ALT_INV_Add0~69_sumout\ <= NOT \Add0~69_sumout\;
\ALT_INV_Add3~77_sumout\ <= NOT \Add3~77_sumout\;
\ALT_INV_Add0~65_sumout\ <= NOT \Add0~65_sumout\;
\ALT_INV_Add3~73_sumout\ <= NOT \Add3~73_sumout\;
\ALT_INV_Add0~61_sumout\ <= NOT \Add0~61_sumout\;
\ALT_INV_Add3~69_sumout\ <= NOT \Add3~69_sumout\;
\ALT_INV_Add0~57_sumout\ <= NOT \Add0~57_sumout\;
\ALT_INV_Add3~65_sumout\ <= NOT \Add3~65_sumout\;
\ALT_INV_Add0~53_sumout\ <= NOT \Add0~53_sumout\;
\ALT_INV_Add3~61_sumout\ <= NOT \Add3~61_sumout\;
\ALT_INV_Add0~49_sumout\ <= NOT \Add0~49_sumout\;
\ALT_INV_Add3~57_sumout\ <= NOT \Add3~57_sumout\;
\ALT_INV_Add0~45_sumout\ <= NOT \Add0~45_sumout\;
\ALT_INV_Add3~53_sumout\ <= NOT \Add3~53_sumout\;
\ALT_INV_Add0~41_sumout\ <= NOT \Add0~41_sumout\;
\ALT_INV_Add3~49_sumout\ <= NOT \Add3~49_sumout\;
\ALT_INV_Add0~37_sumout\ <= NOT \Add0~37_sumout\;
\ALT_INV_Add3~45_sumout\ <= NOT \Add3~45_sumout\;
\ALT_INV_Add0~33_sumout\ <= NOT \Add0~33_sumout\;
\ALT_INV_Add3~41_sumout\ <= NOT \Add3~41_sumout\;
\ALT_INV_Add0~29_sumout\ <= NOT \Add0~29_sumout\;
\ALT_INV_Add3~37_sumout\ <= NOT \Add3~37_sumout\;
\ALT_INV_Add0~25_sumout\ <= NOT \Add0~25_sumout\;
\ALT_INV_Add3~33_sumout\ <= NOT \Add3~33_sumout\;
\ALT_INV_Add0~21_sumout\ <= NOT \Add0~21_sumout\;
\ALT_INV_Add3~29_sumout\ <= NOT \Add3~29_sumout\;
\ALT_INV_Add0~17_sumout\ <= NOT \Add0~17_sumout\;
\ALT_INV_Add3~25_sumout\ <= NOT \Add3~25_sumout\;
\ALT_INV_Add0~13_sumout\ <= NOT \Add0~13_sumout\;
\ALT_INV_Add3~21_sumout\ <= NOT \Add3~21_sumout\;
\ALT_INV_Add0~9_sumout\ <= NOT \Add0~9_sumout\;
\ALT_INV_Add3~17_sumout\ <= NOT \Add3~17_sumout\;
\ALT_INV_Add0~5_sumout\ <= NOT \Add0~5_sumout\;
\ALT_INV_Add3~13_sumout\ <= NOT \Add3~13_sumout\;
\ALT_INV_R.incPC~q\ <= NOT \R.incPC~q\;
\ALT_INV_Add0~1_sumout\ <= NOT \Add0~1_sumout\;
\ALT_INV_Add3~9_sumout\ <= NOT \Add3~9_sumout\;
\ALT_INV_ShiftRight0~7_OTERM233DUPLICATE_q\ <= NOT \ShiftRight0~7_OTERM233DUPLICATE_q\;
\ALT_INV_RegFile[16][23]~DUPLICATE_q\ <= NOT \RegFile[16][23]~DUPLICATE_q\;
\ALT_INV_RegFile[18][20]~DUPLICATE_q\ <= NOT \RegFile[18][20]~DUPLICATE_q\;
\ALT_INV_RegFile[10][18]~DUPLICATE_q\ <= NOT \RegFile[10][18]~DUPLICATE_q\;
\ALT_INV_RegFile[18][31]~DUPLICATE_q\ <= NOT \RegFile[18][31]~DUPLICATE_q\;
\ALT_INV_RegFile[16][5]~DUPLICATE_q\ <= NOT \RegFile[16][5]~DUPLICATE_q\;
\ALT_INV_RegFile[11][11]~DUPLICATE_q\ <= NOT \RegFile[11][11]~DUPLICATE_q\;
\ALT_INV_RegFile[26][27]~DUPLICATE_q\ <= NOT \RegFile[26][27]~DUPLICATE_q\;
\ALT_INV_RegFile[10][10]~DUPLICATE_q\ <= NOT \RegFile[10][10]~DUPLICATE_q\;
\ALT_INV_RegFile[10][26]~DUPLICATE_q\ <= NOT \RegFile[10][26]~DUPLICATE_q\;
\ALT_INV_RegFile[17][9]~DUPLICATE_q\ <= NOT \RegFile[17][9]~DUPLICATE_q\;
\ALT_INV_RegFile[18][0]~DUPLICATE_q\ <= NOT \RegFile[18][0]~DUPLICATE_q\;
\ALT_INV_RegFile[18][8]~DUPLICATE_q\ <= NOT \RegFile[18][8]~DUPLICATE_q\;
\ALT_INV_RegFile[11][8]~DUPLICATE_q\ <= NOT \RegFile[11][8]~DUPLICATE_q\;
\ALT_INV_RegFile[14][20]~DUPLICATE_q\ <= NOT \RegFile[14][20]~DUPLICATE_q\;
\ALT_INV_RegFile[30][18]~DUPLICATE_q\ <= NOT \RegFile[30][18]~DUPLICATE_q\;
\ALT_INV_RegFile[20][16]~DUPLICATE_q\ <= NOT \RegFile[20][16]~DUPLICATE_q\;
\ALT_INV_RegFile[14][16]~DUPLICATE_q\ <= NOT \RegFile[14][16]~DUPLICATE_q\;
\ALT_INV_RegFile[12][16]~DUPLICATE_q\ <= NOT \RegFile[12][16]~DUPLICATE_q\;
\ALT_INV_RegFile[30][7]~DUPLICATE_q\ <= NOT \RegFile[30][7]~DUPLICATE_q\;
\ALT_INV_RegFile[14][6]~DUPLICATE_q\ <= NOT \RegFile[14][6]~DUPLICATE_q\;
\ALT_INV_RegFile[30][30]~DUPLICATE_q\ <= NOT \RegFile[30][30]~DUPLICATE_q\;
\ALT_INV_RegFile[14][2]~DUPLICATE_q\ <= NOT \RegFile[14][2]~DUPLICATE_q\;
\ALT_INV_RegFile[12][10]~DUPLICATE_q\ <= NOT \RegFile[12][10]~DUPLICATE_q\;
\ALT_INV_RegFile[12][1]~DUPLICATE_q\ <= NOT \RegFile[12][1]~DUPLICATE_q\;
\ALT_INV_RegFile[22][9]~DUPLICATE_q\ <= NOT \RegFile[22][9]~DUPLICATE_q\;
\ALT_INV_RegFile[14][9]~DUPLICATE_q\ <= NOT \RegFile[14][9]~DUPLICATE_q\;
\ALT_INV_RegFile[28][0]~DUPLICATE_q\ <= NOT \RegFile[28][0]~DUPLICATE_q\;
\ALT_INV_RegFile[12][0]~DUPLICATE_q\ <= NOT \RegFile[12][0]~DUPLICATE_q\;
\ALT_INV_RegFile[31][8]~DUPLICATE_q\ <= NOT \RegFile[31][8]~DUPLICATE_q\;
\ALT_INV_R.ctrlState.DataAccess0~DUPLICATE_q\ <= NOT \R.ctrlState.DataAccess0~DUPLICATE_q\;
\ALT_INV_RegFile[1][20]~DUPLICATE_q\ <= NOT \RegFile[1][20]~DUPLICATE_q\;
\ALT_INV_RegFile[1][19]~DUPLICATE_q\ <= NOT \RegFile[1][19]~DUPLICATE_q\;
\ALT_INV_RegFile[6][18]~DUPLICATE_q\ <= NOT \RegFile[6][18]~DUPLICATE_q\;
\ALT_INV_RegFile[4][18]~DUPLICATE_q\ <= NOT \RegFile[4][18]~DUPLICATE_q\;
\ALT_INV_RegFile[1][17]~DUPLICATE_q\ <= NOT \RegFile[1][17]~DUPLICATE_q\;
\ALT_INV_RegFile[5][16]~DUPLICATE_q\ <= NOT \RegFile[5][16]~DUPLICATE_q\;
\ALT_INV_RegFile[2][7]~DUPLICATE_q\ <= NOT \RegFile[2][7]~DUPLICATE_q\;
\ALT_INV_RegFile[6][15]~DUPLICATE_q\ <= NOT \RegFile[6][15]~DUPLICATE_q\;
\ALT_INV_RegFile[1][14]~DUPLICATE_q\ <= NOT \RegFile[1][14]~DUPLICATE_q\;
\ALT_INV_RegFile[1][29]~DUPLICATE_q\ <= NOT \RegFile[1][29]~DUPLICATE_q\;
\ALT_INV_RegFile[2][12]~DUPLICATE_q\ <= NOT \RegFile[2][12]~DUPLICATE_q\;
\ALT_INV_RegFile[6][28]~DUPLICATE_q\ <= NOT \RegFile[6][28]~DUPLICATE_q\;
\ALT_INV_RegFile[2][26]~DUPLICATE_q\ <= NOT \RegFile[2][26]~DUPLICATE_q\;
\ALT_INV_RegFile[7][26]~DUPLICATE_q\ <= NOT \RegFile[7][26]~DUPLICATE_q\;
\ALT_INV_RegFile[6][8]~DUPLICATE_q\ <= NOT \RegFile[6][8]~DUPLICATE_q\;
\ALT_INV_R.aluRes[30]~DUPLICATE_q\ <= NOT \R.aluRes[30]~DUPLICATE_q\;
\ALT_INV_R.aluRes[27]~DUPLICATE_q\ <= NOT \R.aluRes[27]~DUPLICATE_q\;
\ALT_INV_R.aluRes[4]~DUPLICATE_q\ <= NOT \R.aluRes[4]~DUPLICATE_q\;
\ALT_INV_R.aluRes[0]~DUPLICATE_q\ <= NOT \R.aluRes[0]~DUPLICATE_q\;
\ALT_INV_R.aluOp.ALUOpAnd~DUPLICATE_q\ <= NOT \R.aluOp.ALUOpAnd~DUPLICATE_q\;
\ALT_INV_R.aluOp.ALUOpXor~DUPLICATE_q\ <= NOT \R.aluOp.ALUOpXor~DUPLICATE_q\;
\ALT_INV_R.aluData2[25]~DUPLICATE_q\ <= NOT \R.aluData2[25]~DUPLICATE_q\;
\ALT_INV_R.aluData2[13]~DUPLICATE_q\ <= NOT \R.aluData2[13]~DUPLICATE_q\;
\ALT_INV_R.curPC[0]~DUPLICATE_q\ <= NOT \R.curPC[0]~DUPLICATE_q\;
\ALT_INV_R.curPC[31]~DUPLICATE_q\ <= NOT \R.curPC[31]~DUPLICATE_q\;
\ALT_INV_R.curPC[30]~DUPLICATE_q\ <= NOT \R.curPC[30]~DUPLICATE_q\;
\ALT_INV_R.curPC[21]~DUPLICATE_q\ <= NOT \R.curPC[21]~DUPLICATE_q\;
\ALT_INV_Comb:vRegWriteData[18]~1_RESYN1740_BDD1741\ <= NOT \Comb:vRegWriteData[18]~1_RESYN1740_BDD1741\;
\ALT_INV_Comb:vRegWriteData[18]~1_RESYN1738_BDD1739\ <= NOT \Comb:vRegWriteData[18]~1_RESYN1738_BDD1739\;
\ALT_INV_Comb:vRegWriteData[18]~1_RESYN1736_BDD1737\ <= NOT \Comb:vRegWriteData[18]~1_RESYN1736_BDD1737\;
\ALT_INV_Comb:vRegWriteData[8]~1_RESYN1734_BDD1735\ <= NOT \Comb:vRegWriteData[8]~1_RESYN1734_BDD1735\;
\ALT_INV_Comb:vRegWriteData[8]~1_RESYN1732_BDD1733\ <= NOT \Comb:vRegWriteData[8]~1_RESYN1732_BDD1733\;
\ALT_INV_Comb:vRegWriteData[8]~1_RESYN1730_BDD1731\ <= NOT \Comb:vRegWriteData[8]~1_RESYN1730_BDD1731\;
\ALT_INV_Comb:vRegWriteData[16]~0_RESYN1728_BDD1729\ <= NOT \Comb:vRegWriteData[16]~0_RESYN1728_BDD1729\;
\ALT_INV_Comb:vRegWriteData[16]~0_RESYN1726_BDD1727\ <= NOT \Comb:vRegWriteData[16]~0_RESYN1726_BDD1727\;
\ALT_INV_Comb:vRegWriteData[16]~0_RESYN1724_BDD1725\ <= NOT \Comb:vRegWriteData[16]~0_RESYN1724_BDD1725\;
\ALT_INV_vAluRes~7_RESYN1076_RESYN1132_BDD1133\ <= NOT \vAluRes~7_RESYN1076_RESYN1132_BDD1133\;
\ALT_INV_Comb:vRegWriteData[21]~1_RESYN1130_BDD1131\ <= NOT \Comb:vRegWriteData[21]~1_RESYN1130_BDD1131\;
\ALT_INV_Comb:vRegWriteData[21]~1_RESYN1128_BDD1129\ <= NOT \Comb:vRegWriteData[21]~1_RESYN1128_BDD1129\;
\ALT_INV_Comb:vRegWriteData[21]~1_RESYN1126_BDD1127\ <= NOT \Comb:vRegWriteData[21]~1_RESYN1126_BDD1127\;
\ALT_INV_Comb:vRegWriteData[17]~1_RESYN1124_BDD1125\ <= NOT \Comb:vRegWriteData[17]~1_RESYN1124_BDD1125\;
\ALT_INV_Comb:vRegWriteData[17]~1_RESYN1122_BDD1123\ <= NOT \Comb:vRegWriteData[17]~1_RESYN1122_BDD1123\;
\ALT_INV_Comb:vRegWriteData[17]~1_RESYN1120_BDD1121\ <= NOT \Comb:vRegWriteData[17]~1_RESYN1120_BDD1121\;
\ALT_INV_Comb:vRegWriteData[7]~0_RESYN1118_BDD1119\ <= NOT \Comb:vRegWriteData[7]~0_RESYN1118_BDD1119\;
\ALT_INV_Selector25~6_RESYN1116_BDD1117\ <= NOT \Selector25~6_RESYN1116_BDD1117\;
\ALT_INV_Comb:vRegWriteData[23]~2_RESYN1114_BDD1115\ <= NOT \Comb:vRegWriteData[23]~2_RESYN1114_BDD1115\;
\ALT_INV_Comb:vRegWriteData[22]~2_RESYN1112_BDD1113\ <= NOT \Comb:vRegWriteData[22]~2_RESYN1112_BDD1113\;
\ALT_INV_Comb:vRegWriteData[20]~2_RESYN1110_BDD1111\ <= NOT \Comb:vRegWriteData[20]~2_RESYN1110_BDD1111\;
\ALT_INV_Comb:vRegWriteData[27]~2_RESYN1108_BDD1109\ <= NOT \Comb:vRegWriteData[27]~2_RESYN1108_BDD1109\;
\ALT_INV_Comb:vRegWriteData[25]~2_RESYN1106_BDD1107\ <= NOT \Comb:vRegWriteData[25]~2_RESYN1106_BDD1107\;
\ALT_INV_Comb:vRegWriteData[24]~3_RESYN1104_BDD1105\ <= NOT \Comb:vRegWriteData[24]~3_RESYN1104_BDD1105\;
\ALT_INV_Equal3~5_RESYN1102_BDD1103\ <= NOT \Equal3~5_RESYN1102_BDD1103\;
\ALT_INV_Equal3~5_RESYN1100_BDD1101\ <= NOT \Equal3~5_RESYN1100_BDD1101\;
\ALT_INV_Comb:vRegWriteData[6]~0_RESYN1098_BDD1099\ <= NOT \Comb:vRegWriteData[6]~0_RESYN1098_BDD1099\;
\ALT_INV_Comb:vRegWriteData[14]~1_RESYN1096_BDD1097\ <= NOT \Comb:vRegWriteData[14]~1_RESYN1096_BDD1097\;
\ALT_INV_Comb:vRegWriteData[14]~1_RESYN1094_BDD1095\ <= NOT \Comb:vRegWriteData[14]~1_RESYN1094_BDD1095\;
\ALT_INV_Comb:vRegWriteData[5]~0_RESYN1092_BDD1093\ <= NOT \Comb:vRegWriteData[5]~0_RESYN1092_BDD1093\;
\ALT_INV_Comb:vRegWriteData[4]~0_RESYN1090_BDD1091\ <= NOT \Comb:vRegWriteData[4]~0_RESYN1090_BDD1091\;
\ALT_INV_Comb:vRegWriteData[12]~1_RESYN1088_BDD1089\ <= NOT \Comb:vRegWriteData[12]~1_RESYN1088_BDD1089\;
\ALT_INV_Comb:vRegWriteData[12]~1_RESYN1086_BDD1087\ <= NOT \Comb:vRegWriteData[12]~1_RESYN1086_BDD1087\;
\ALT_INV_Comb:vRegWriteData[3]~0_RESYN1084_BDD1085\ <= NOT \Comb:vRegWriteData[3]~0_RESYN1084_BDD1085\;
\ALT_INV_Comb:vRegWriteData[2]~0_RESYN1082_BDD1083\ <= NOT \Comb:vRegWriteData[2]~0_RESYN1082_BDD1083\;
\ALT_INV_Comb:vRegWriteData[9]~1_RESYN1080_BDD1081\ <= NOT \Comb:vRegWriteData[9]~1_RESYN1080_BDD1081\;
\ALT_INV_Comb:vRegWriteData[9]~1_RESYN1078_BDD1079\ <= NOT \Comb:vRegWriteData[9]~1_RESYN1078_BDD1079\;
\ALT_INV_vAluRes~7_RESYN1076_BDD1077\ <= NOT \vAluRes~7_RESYN1076_BDD1077\;
\ALT_INV_vAluRes~6_RESYN1072_BDD1073\ <= NOT \vAluRes~6_RESYN1072_BDD1073\;
\ALT_INV_vAluRes~5_RESYN1070_BDD1071\ <= NOT \vAluRes~5_RESYN1070_BDD1071\;
\ALT_INV_vAluRes~4_RESYN1068_BDD1069\ <= NOT \vAluRes~4_RESYN1068_BDD1069\;
\ALT_INV_vAluRes~3_RESYN1066_BDD1067\ <= NOT \vAluRes~3_RESYN1066_BDD1067\;
\ALT_INV_vAluRes~2_RESYN1064_BDD1065\ <= NOT \vAluRes~2_RESYN1064_BDD1065\;
\ALT_INV_vAluRes~1_RESYN1062_BDD1063\ <= NOT \vAluRes~1_RESYN1062_BDD1063\;
\ALT_INV_Selector32~7_RESYN1060_BDD1061\ <= NOT \Selector32~7_RESYN1060_BDD1061\;
\ALT_INV_Selector32~7_RESYN1058_BDD1059\ <= NOT \Selector32~7_RESYN1058_BDD1059\;
\ALT_INV_Selector32~7_RESYN1056_BDD1057\ <= NOT \Selector32~7_RESYN1056_BDD1057\;
\ALT_INV_Equal3~12_RESYN1054_BDD1055\ <= NOT \Equal3~12_RESYN1054_BDD1055\;
\ALT_INV_Comb:vRegWriteData[15]~1_RESYN1048_BDD1049\ <= NOT \Comb:vRegWriteData[15]~1_RESYN1048_BDD1049\;
\ALT_INV_Comb:vRegWriteData[15]~1_RESYN1046_BDD1047\ <= NOT \Comb:vRegWriteData[15]~1_RESYN1046_BDD1047\;
\ALT_INV_Comb:vRegWriteData[13]~1_RESYN1044_BDD1045\ <= NOT \Comb:vRegWriteData[13]~1_RESYN1044_BDD1045\;
\ALT_INV_Comb:vRegWriteData[13]~1_RESYN1042_BDD1043\ <= NOT \Comb:vRegWriteData[13]~1_RESYN1042_BDD1043\;
\ALT_INV_Comb:vRegWriteData[11]~1_RESYN1040_BDD1041\ <= NOT \Comb:vRegWriteData[11]~1_RESYN1040_BDD1041\;
\ALT_INV_Comb:vRegWriteData[11]~1_RESYN1038_BDD1039\ <= NOT \Comb:vRegWriteData[11]~1_RESYN1038_BDD1039\;
\ALT_INV_Comb:vJumpAdr[30]~0_RESYN1036_BDD1037\ <= NOT \Comb:vJumpAdr[30]~0_RESYN1036_BDD1037\;
\ALT_INV_Comb:vJumpAdr[29]~0_RESYN1034_BDD1035\ <= NOT \Comb:vJumpAdr[29]~0_RESYN1034_BDD1035\;
\ALT_INV_Comb:vJumpAdr[28]~0_RESYN1032_BDD1033\ <= NOT \Comb:vJumpAdr[28]~0_RESYN1032_BDD1033\;
\ALT_INV_Comb:vJumpAdr[27]~0_RESYN1030_BDD1031\ <= NOT \Comb:vJumpAdr[27]~0_RESYN1030_BDD1031\;
\ALT_INV_Comb:vJumpAdr[22]~0_RESYN1028_BDD1029\ <= NOT \Comb:vJumpAdr[22]~0_RESYN1028_BDD1029\;
\ALT_INV_Add2~17_OTERM727_OTERM841\ <= NOT \Add2~17_OTERM727_OTERM841\;
\ALT_INV_Add2~1_OTERM735_OTERM839\ <= NOT \Add2~1_OTERM735_OTERM839\;
\ALT_INV_Add2~1_OTERM735_OTERM837\ <= NOT \Add2~1_OTERM735_OTERM837\;
\ALT_INV_Add2~25_OTERM723_OTERM835\ <= NOT \Add2~25_OTERM723_OTERM835\;
\ALT_INV_Add2~25_OTERM723_OTERM833\ <= NOT \Add2~25_OTERM723_OTERM833\;
\ALT_INV_Add2~25_OTERM723_OTERM831\ <= NOT \Add2~25_OTERM723_OTERM831\;
\ALT_INV_Add2~25_OTERM723_OTERM829\ <= NOT \Add2~25_OTERM723_OTERM829\;
\ALT_INV_Add2~33_OTERM719_OTERM827\ <= NOT \Add2~33_OTERM719_OTERM827\;
\ALT_INV_Add2~33_OTERM719_OTERM825\ <= NOT \Add2~33_OTERM719_OTERM825\;
\ALT_INV_Add2~33_OTERM719_OTERM823\ <= NOT \Add2~33_OTERM719_OTERM823\;
\ALT_INV_Add2~33_OTERM719_OTERM821\ <= NOT \Add2~33_OTERM719_OTERM821\;
\ALT_INV_Add2~41_OTERM715_OTERM819\ <= NOT \Add2~41_OTERM715_OTERM819\;
\ALT_INV_Add2~41_OTERM715_OTERM817\ <= NOT \Add2~41_OTERM715_OTERM817\;
\ALT_INV_Add2~57_OTERM707_OTERM815\ <= NOT \Add2~57_OTERM707_OTERM815\;
\ALT_INV_Add2~57_OTERM707_OTERM813\ <= NOT \Add2~57_OTERM707_OTERM813\;
\ALT_INV_Add2~65_OTERM703_OTERM811\ <= NOT \Add2~65_OTERM703_OTERM811\;
\ALT_INV_Add2~65_OTERM703_OTERM809\ <= NOT \Add2~65_OTERM703_OTERM809\;
\ALT_INV_Add2~65_OTERM703_OTERM807\ <= NOT \Add2~65_OTERM703_OTERM807\;
\ALT_INV_Add2~65_OTERM703_OTERM805\ <= NOT \Add2~65_OTERM703_OTERM805\;
\ALT_INV_Selector19~1_OTERM751_OTERM803\ <= NOT \Selector19~1_OTERM751_OTERM803\;
\ALT_INV_Selector25~3_OTERM797\ <= NOT \Selector25~3_OTERM797\;
\ALT_INV_Selector16~1_OTERM793\ <= NOT \Selector16~1_OTERM793\;
\ALT_INV_ShiftLeft0~12_OTERM791\ <= NOT \ShiftLeft0~12_OTERM791\;
\ALT_INV_ShiftLeft0~38_OTERM789\ <= NOT \ShiftLeft0~38_OTERM789\;
\ALT_INV_Selector1~0_OTERM771\ <= NOT \Selector1~0_OTERM771\;
\ALT_INV_Selector20~0_OTERM769\ <= NOT \Selector20~0_OTERM769\;
\ALT_INV_ShiftLeft0~55_OTERM767\ <= NOT \ShiftLeft0~55_OTERM767\;
\ALT_INV_ShiftLeft0~53_OTERM765\ <= NOT \ShiftLeft0~53_OTERM765\;
\ALT_INV_ShiftLeft0~51_OTERM763\ <= NOT \ShiftLeft0~51_OTERM763\;
\ALT_INV_ShiftLeft0~49_OTERM761\ <= NOT \ShiftLeft0~49_OTERM761\;
\ALT_INV_ShiftLeft0~47_OTERM759\ <= NOT \ShiftLeft0~47_OTERM759\;
\ALT_INV_ShiftLeft0~45_OTERM757\ <= NOT \ShiftLeft0~45_OTERM757\;
\ALT_INV_ShiftLeft0~40_OTERM755\ <= NOT \ShiftLeft0~40_OTERM755\;
\ALT_INV_ShiftLeft0~14_OTERM753\ <= NOT \ShiftLeft0~14_OTERM753\;
\ALT_INV_Selector22~0_OTERM475_OTERM749\ <= NOT \Selector22~0_OTERM475_OTERM749\;
\ALT_INV_Selector22~0_OTERM475_OTERM747\ <= NOT \Selector22~0_OTERM475_OTERM747\;
\ALT_INV_ShiftRight1~38_OTERM439_OTERM745\ <= NOT \ShiftRight1~38_OTERM439_OTERM745\;
\ALT_INV_Selector15~2_OTERM741\ <= NOT \Selector15~2_OTERM741\;
\ALT_INV_ShiftLeft0~26_OTERM739\ <= NOT \ShiftLeft0~26_OTERM739\;
\ALT_INV_ShiftLeft0~22_OTERM737\ <= NOT \ShiftLeft0~22_OTERM737\;
\ALT_INV_ShiftLeft0~36_OTERM603\ <= NOT \ShiftLeft0~36_OTERM603\;
\ALT_INV_ShiftLeft0~30_OTERM601\ <= NOT \ShiftLeft0~30_OTERM601\;
\ALT_INV_Selector31~5_OTERM599\ <= NOT \Selector31~5_OTERM599\;
\ALT_INV_R.statusReg[0]_OTERM11_OTERM377_OTERM597\ <= NOT \R.statusReg[0]_OTERM11_OTERM377_OTERM597\;
\ALT_INV_R.statusReg[0]_OTERM11_OTERM377_OTERM595\ <= NOT \R.statusReg[0]_OTERM11_OTERM377_OTERM595\;
\ALT_INV_R.statusReg[0]_OTERM11_OTERM377_OTERM593\ <= NOT \R.statusReg[0]_OTERM11_OTERM377_OTERM593\;
\ALT_INV_Selector31~0_NEW_REG348_OTERM569\ <= NOT \Selector31~0_NEW_REG348_OTERM569\;
\ALT_INV_R.statusReg[0]_OTERM7_OTERM491\ <= NOT \R.statusReg[0]_OTERM7_OTERM491\;
\ALT_INV_R.statusReg[0]_OTERM7_OTERM489\ <= NOT \R.statusReg[0]_OTERM7_OTERM489\;
\ALT_INV_R.statusReg[0]_OTERM7_OTERM487\ <= NOT \R.statusReg[0]_OTERM7_OTERM487\;
\ALT_INV_R.statusReg[0]_OTERM7_OTERM485\ <= NOT \R.statusReg[0]_OTERM7_OTERM485\;
\ALT_INV_R.statusReg[0]_OTERM7_OTERM483\ <= NOT \R.statusReg[0]_OTERM7_OTERM483\;
\ALT_INV_R.statusReg[0]_OTERM7_OTERM481\ <= NOT \R.statusReg[0]_OTERM7_OTERM481\;
\ALT_INV_Selector22~0_RTM0477_combout\ <= NOT \Selector22~0_RTM0477_combout\;
\ALT_INV_R.statusReg[0]_OTERM9_OTERM473\ <= NOT \R.statusReg[0]_OTERM9_OTERM473\;
\ALT_INV_R.statusReg[0]_OTERM9_OTERM471\ <= NOT \R.statusReg[0]_OTERM9_OTERM471\;
\ALT_INV_R.statusReg[0]_OTERM9_OTERM469\ <= NOT \R.statusReg[0]_OTERM9_OTERM469\;
\ALT_INV_R.statusReg[0]_OTERM9_OTERM467\ <= NOT \R.statusReg[0]_OTERM9_OTERM467\;
\ALT_INV_R.statusReg[0]_OTERM9_OTERM465\ <= NOT \R.statusReg[0]_OTERM9_OTERM465\;
\ALT_INV_R.statusReg[0]_OTERM9_OTERM463\ <= NOT \R.statusReg[0]_OTERM9_OTERM463\;
\ALT_INV_ShiftLeft0~9_OTERM461\ <= NOT \ShiftLeft0~9_OTERM461\;
\ALT_INV_Selector18~1_OTERM431\ <= NOT \Selector18~1_OTERM431\;
\ALT_INV_Selector22~1_OTERM427\ <= NOT \Selector22~1_OTERM427\;
\ALT_INV_Selector23~3_OTERM423\ <= NOT \Selector23~3_OTERM423\;
\ALT_INV_Selector24~0_OTERM419\ <= NOT \Selector24~0_OTERM419\;
\ALT_INV_Selector26~2_OTERM415\ <= NOT \Selector26~2_OTERM415\;
\ALT_INV_Selector27~2_OTERM411\ <= NOT \Selector27~2_OTERM411\;
\ALT_INV_Selector29~0_OTERM407\ <= NOT \Selector29~0_OTERM407\;
\ALT_INV_Selector30~1_OTERM403\ <= NOT \Selector30~1_OTERM403\;
\ALT_INV_Selector31~2_OTERM399\ <= NOT \Selector31~2_OTERM399\;
\ALT_INV_Selector32~4_OTERM397\ <= NOT \Selector32~4_OTERM397\;
\ALT_INV_Selector12~2_OTERM395\ <= NOT \Selector12~2_OTERM395\;
\ALT_INV_Selector16~0_OTERM393\ <= NOT \Selector16~0_OTERM393\;
\ALT_INV_Selector17~0_OTERM391\ <= NOT \Selector17~0_OTERM391\;
\ALT_INV_Selector28~1_OTERM387\ <= NOT \Selector28~1_OTERM387\;
\ALT_INV_Selector27~0_OTERM385\ <= NOT \Selector27~0_OTERM385\;
\ALT_INV_Selector31~7_OTERM383\ <= NOT \Selector31~7_OTERM383\;
\ALT_INV_Selector31~6_OTERM381\ <= NOT \Selector31~6_OTERM381\;
\ALT_INV_Selector32~3_OTERM379\ <= NOT \Selector32~3_OTERM379\;
\ALT_INV_R.statusReg[0]_OTERM11_OTERM375\ <= NOT \R.statusReg[0]_OTERM11_OTERM375\;
\ALT_INV_R.statusReg[0]_OTERM11_OTERM373\ <= NOT \R.statusReg[0]_OTERM11_OTERM373\;
\ALT_INV_R.statusReg[0]_OTERM11_OTERM371\ <= NOT \R.statusReg[0]_OTERM11_OTERM371\;
\ALT_INV_R.statusReg[0]_OTERM11_OTERM369\ <= NOT \R.statusReg[0]_OTERM11_OTERM369\;
\ALT_INV_R.statusReg[0]_OTERM11_OTERM367\ <= NOT \R.statusReg[0]_OTERM11_OTERM367\;
\ALT_INV_R.aluOp.ALUOpSRA_OTERM363\ <= NOT \R.aluOp.ALUOpSRA_OTERM363\;
\ALT_INV_R.aluOp.ALUOpSRL_OTERM361\ <= NOT \R.aluOp.ALUOpSRL_OTERM361\;
\ALT_INV_R.aluOp.ALUOpSLL_OTERM359\ <= NOT \R.aluOp.ALUOpSLL_OTERM359\;
\ALT_INV_R.aluOp.ALUOpAnd_OTERM357\ <= NOT \R.aluOp.ALUOpAnd_OTERM357\;
\ALT_INV_R.aluOp.ALUOpXor_OTERM355\ <= NOT \R.aluOp.ALUOpXor_OTERM355\;
\ALT_INV_R.aluOp.ALUOpOr_OTERM353\ <= NOT \R.aluOp.ALUOpOr_OTERM353\;
\ALT_INV_Selector31~0_OTERM349\ <= NOT \Selector31~0_OTERM349\;
\ALT_INV_LessThan1~22_OTERM347\ <= NOT \LessThan1~22_OTERM347\;
\ALT_INV_LessThan1~0_OTERM343\ <= NOT \LessThan1~0_OTERM343\;
\ALT_INV_LessThan1~20_OTERM341\ <= NOT \LessThan1~20_OTERM341\;
\ALT_INV_LessThan1~1_OTERM337\ <= NOT \LessThan1~1_OTERM337\;
\ALT_INV_LessThan1~21_OTERM335\ <= NOT \LessThan1~21_OTERM335\;
\ALT_INV_LessThan1~2_OTERM331\ <= NOT \LessThan1~2_OTERM331\;
\ALT_INV_LessThan1~24_OTERM329\ <= NOT \LessThan1~24_OTERM329\;
\ALT_INV_LessThan1~3_OTERM325\ <= NOT \LessThan1~3_OTERM325\;
\ALT_INV_LessThan1~18_OTERM321\ <= NOT \LessThan1~18_OTERM321\;
\ALT_INV_LessThan1~4_OTERM319\ <= NOT \LessThan1~4_OTERM319\;
\ALT_INV_LessThan1~25_OTERM317\ <= NOT \LessThan1~25_OTERM317\;
\ALT_INV_LessThan1~5_OTERM313\ <= NOT \LessThan1~5_OTERM313\;
\ALT_INV_LessThan1~16_OTERM311\ <= NOT \LessThan1~16_OTERM311\;
\ALT_INV_LessThan1~7_OTERM307\ <= NOT \LessThan1~7_OTERM307\;
\ALT_INV_LessThan1~14_OTERM305\ <= NOT \LessThan1~14_OTERM305\;
\ALT_INV_LessThan1~8_OTERM301\ <= NOT \LessThan1~8_OTERM301\;
\ALT_INV_ShiftLeft0~34_OTERM299\ <= NOT \ShiftLeft0~34_OTERM299\;
\ALT_INV_ShiftLeft0~32_OTERM297\ <= NOT \ShiftLeft0~32_OTERM297\;
\ALT_INV_ShiftLeft0~28_OTERM295\ <= NOT \ShiftLeft0~28_OTERM295\;
\ALT_INV_ShiftLeft0~24_OTERM293\ <= NOT \ShiftLeft0~24_OTERM293\;
\ALT_INV_ShiftLeft0~20_OTERM291\ <= NOT \ShiftLeft0~20_OTERM291\;
\ALT_INV_ShiftLeft0~18_OTERM289\ <= NOT \ShiftLeft0~18_OTERM289\;
\ALT_INV_ShiftLeft0~16_OTERM287\ <= NOT \ShiftLeft0~16_OTERM287\;
\ALT_INV_ShiftLeft0~13_OTERM285\ <= NOT \ShiftLeft0~13_OTERM285\;
\ALT_INV_ShiftRight1~37_OTERM283\ <= NOT \ShiftRight1~37_OTERM283\;
\ALT_INV_ShiftRight1~36_OTERM281\ <= NOT \ShiftRight1~36_OTERM281\;
\ALT_INV_ShiftRight1~35_OTERM279\ <= NOT \ShiftRight1~35_OTERM279\;
\ALT_INV_ShiftRight1~25_OTERM277\ <= NOT \ShiftRight1~25_OTERM277\;
\ALT_INV_ShiftRight1~23_OTERM275\ <= NOT \ShiftRight1~23_OTERM275\;
\ALT_INV_ShiftRight1~22_OTERM273\ <= NOT \ShiftRight1~22_OTERM273\;
\ALT_INV_ShiftRight1~21_OTERM271\ <= NOT \ShiftRight1~21_OTERM271\;
\ALT_INV_ShiftRight1~18_OTERM269\ <= NOT \ShiftRight1~18_OTERM269\;
\ALT_INV_ShiftRight1~17_OTERM267\ <= NOT \ShiftRight1~17_OTERM267\;
\ALT_INV_ShiftRight1~10_OTERM265\ <= NOT \ShiftRight1~10_OTERM265\;
\ALT_INV_ShiftLeft0~0_OTERM263\ <= NOT \ShiftLeft0~0_OTERM263\;
\ALT_INV_ShiftRight1~8_OTERM261\ <= NOT \ShiftRight1~8_OTERM261\;
\ALT_INV_ShiftRight1~7_OTERM259\ <= NOT \ShiftRight1~7_OTERM259\;
\ALT_INV_ShiftRight1~0_OTERM257\ <= NOT \ShiftRight1~0_OTERM257\;
\ALT_INV_ShiftLeft0~1_OTERM255\ <= NOT \ShiftLeft0~1_OTERM255\;
\ALT_INV_LessThan1~9_OTERM253\ <= NOT \LessThan1~9_OTERM253\;
\ALT_INV_ShiftLeft0~6_OTERM243\ <= NOT \ShiftLeft0~6_OTERM243\;
\ALT_INV_ShiftLeft0~4_OTERM237\ <= NOT \ShiftLeft0~4_OTERM237\;
\ALT_INV_ShiftRight0~7_OTERM233\ <= NOT \ShiftRight0~7_OTERM233\;
\ALT_INV_ShiftLeft0~3_OTERM223\ <= NOT \ShiftLeft0~3_OTERM223\;
\ALT_INV_ShiftLeft0~2_OTERM221\ <= NOT \ShiftLeft0~2_OTERM221\;
\ALT_INV_ShiftRight1~5_OTERM219\ <= NOT \ShiftRight1~5_OTERM219\;
\ALT_INV_LessThan1~11_OTERM217\ <= NOT \LessThan1~11_OTERM217\;
\ALT_INV_LessThan1~10_OTERM213\ <= NOT \LessThan1~10_OTERM213\;
\ALT_INV_ShiftLeft0~10_OTERM211\ <= NOT \ShiftLeft0~10_OTERM211\;
\ALT_INV_ShiftRight1~16_OTERM209\ <= NOT \ShiftRight1~16_OTERM209\;
\ALT_INV_ShiftLeft0~8_OTERM207\ <= NOT \ShiftLeft0~8_OTERM207\;
\ALT_INV_ShiftLeft0~7_OTERM205\ <= NOT \ShiftLeft0~7_OTERM205\;
\ALT_INV_ShiftLeft0~5_OTERM203\ <= NOT \ShiftLeft0~5_OTERM203\;
\ALT_INV_ShiftRight1~15_OTERM199\ <= NOT \ShiftRight1~15_OTERM199\;
\ALT_INV_ShiftRight1~6_OTERM197\ <= NOT \ShiftRight1~6_OTERM197\;
\ALT_INV_LessThan1~15_OTERM195\ <= NOT \LessThan1~15_OTERM195\;
\ALT_INV_LessThan1~12_OTERM191\ <= NOT \LessThan1~12_OTERM191\;
\ALT_INV_ShiftRight1~12_OTERM57\ <= NOT \ShiftRight1~12_OTERM57\;
\ALT_INV_LessThan1~34_OTERM55\ <= NOT \LessThan1~34_OTERM55\;
\ALT_INV_LessThan1~28_OTERM51\ <= NOT \LessThan1~28_OTERM51\;
\ALT_INV_ShiftRight1~2_OTERM49\ <= NOT \ShiftRight1~2_OTERM49\;
\ALT_INV_LessThan1~29_OTERM47\ <= NOT \LessThan1~29_OTERM47\;
\ALT_INV_ShiftRight1~31_OTERM45\ <= NOT \ShiftRight1~31_OTERM45\;
\ALT_INV_LessThan1~30_OTERM43\ <= NOT \LessThan1~30_OTERM43\;
\ALT_INV_ShiftLeft0~42_OTERM41\ <= NOT \ShiftLeft0~42_OTERM41\;
\ALT_INV_ShiftRight1~30_OTERM39\ <= NOT \ShiftRight1~30_OTERM39\;
\ALT_INV_ShiftRight1~26_OTERM37\ <= NOT \ShiftRight1~26_OTERM37\;
\ALT_INV_ShiftRight1~11_OTERM35\ <= NOT \ShiftRight1~11_OTERM35\;
\ALT_INV_ShiftRight1~1_OTERM33\ <= NOT \ShiftRight1~1_OTERM33\;
\ALT_INV_ShiftRight0~4_OTERM31\ <= NOT \ShiftRight0~4_OTERM31\;
\ALT_INV_ShiftRight0~2_OTERM25\ <= NOT \ShiftRight0~2_OTERM25\;
\ALT_INV_ShiftRight1~28_OTERM23\ <= NOT \ShiftRight1~28_OTERM23\;
\ALT_INV_ShiftRight1~32_OTERM21\ <= NOT \ShiftRight1~32_OTERM21\;
\ALT_INV_ShiftRight1~27_OTERM19\ <= NOT \ShiftRight1~27_OTERM19\;
\ALT_INV_ShiftRight0~0_OTERM17\ <= NOT \ShiftRight0~0_OTERM17\;
\ALT_INV_ShiftRight1~13_OTERM15\ <= NOT \ShiftRight1~13_OTERM15\;
\ALT_INV_ShiftRight1~3_OTERM13\ <= NOT \ShiftRight1~3_OTERM13\;
\ALT_INV_R.statusReg[0]_OTERM5\ <= NOT \R.statusReg[0]_OTERM5\;
\ALT_INV_R.statusReg[0]_OTERM3\ <= NOT \R.statusReg[0]_OTERM3\;
\ALT_INV_R.statusReg[0]_OTERM1\ <= NOT \R.statusReg[0]_OTERM1\;
\ALT_INV_avm_d_readdata[15]~input_o\ <= NOT \avm_d_readdata[15]~input_o\;
\ALT_INV_avm_d_readdata[14]~input_o\ <= NOT \avm_d_readdata[14]~input_o\;
\ALT_INV_avm_d_readdata[13]~input_o\ <= NOT \avm_d_readdata[13]~input_o\;
\ALT_INV_avm_d_readdata[12]~input_o\ <= NOT \avm_d_readdata[12]~input_o\;
\ALT_INV_avm_d_readdata[11]~input_o\ <= NOT \avm_d_readdata[11]~input_o\;
\ALT_INV_avm_d_readdata[10]~input_o\ <= NOT \avm_d_readdata[10]~input_o\;
\ALT_INV_avm_d_readdata[9]~input_o\ <= NOT \avm_d_readdata[9]~input_o\;
\ALT_INV_avm_d_readdata[8]~input_o\ <= NOT \avm_d_readdata[8]~input_o\;
\ALT_INV_avm_d_readdata[7]~input_o\ <= NOT \avm_d_readdata[7]~input_o\;
\ALT_INV_avm_d_readdata[30]~input_o\ <= NOT \avm_d_readdata[30]~input_o\;
\ALT_INV_avm_d_readdata[22]~input_o\ <= NOT \avm_d_readdata[22]~input_o\;
\ALT_INV_avm_d_readdata[6]~input_o\ <= NOT \avm_d_readdata[6]~input_o\;
\ALT_INV_avm_d_readdata[29]~input_o\ <= NOT \avm_d_readdata[29]~input_o\;
\ALT_INV_avm_d_readdata[21]~input_o\ <= NOT \avm_d_readdata[21]~input_o\;
\ALT_INV_avm_d_readdata[5]~input_o\ <= NOT \avm_d_readdata[5]~input_o\;
\ALT_INV_avm_d_readdata[28]~input_o\ <= NOT \avm_d_readdata[28]~input_o\;
\ALT_INV_avm_d_readdata[20]~input_o\ <= NOT \avm_d_readdata[20]~input_o\;
\ALT_INV_avm_d_readdata[4]~input_o\ <= NOT \avm_d_readdata[4]~input_o\;
\ALT_INV_avm_d_readdata[27]~input_o\ <= NOT \avm_d_readdata[27]~input_o\;
\ALT_INV_avm_d_readdata[19]~input_o\ <= NOT \avm_d_readdata[19]~input_o\;
\ALT_INV_avm_d_readdata[3]~input_o\ <= NOT \avm_d_readdata[3]~input_o\;
\ALT_INV_avm_d_readdata[26]~input_o\ <= NOT \avm_d_readdata[26]~input_o\;
\ALT_INV_avm_d_readdata[18]~input_o\ <= NOT \avm_d_readdata[18]~input_o\;
\ALT_INV_avm_d_readdata[2]~input_o\ <= NOT \avm_d_readdata[2]~input_o\;
\ALT_INV_avm_d_readdata[25]~input_o\ <= NOT \avm_d_readdata[25]~input_o\;
\ALT_INV_avm_d_readdata[17]~input_o\ <= NOT \avm_d_readdata[17]~input_o\;
\ALT_INV_avm_d_readdata[1]~input_o\ <= NOT \avm_d_readdata[1]~input_o\;
\ALT_INV_avm_d_readdata[24]~input_o\ <= NOT \avm_d_readdata[24]~input_o\;
\ALT_INV_avm_d_readdata[16]~input_o\ <= NOT \avm_d_readdata[16]~input_o\;
\ALT_INV_avm_d_readdata[23]~input_o\ <= NOT \avm_d_readdata[23]~input_o\;
\ALT_INV_avm_d_readdata[31]~input_o\ <= NOT \avm_d_readdata[31]~input_o\;
\ALT_INV_avm_d_readdata[0]~input_o\ <= NOT \avm_d_readdata[0]~input_o\;
\ALT_INV_Equal3~15_combout\ <= NOT \Equal3~15_combout\;
\ALT_INV_Equal3~14_combout\ <= NOT \Equal3~14_combout\;
\ALT_INV_Comb:vRegWriteData[23]~3_combout\ <= NOT \Comb:vRegWriteData[23]~3_combout\;
\ALT_INV_Comb:vRegWriteData[23]~2_combout\ <= NOT \Comb:vRegWriteData[23]~2_combout\;
\ALT_INV_Comb:vRegWriteData[23]~1_combout\ <= NOT \Comb:vRegWriteData[23]~1_combout\;
\ALT_INV_Comb:vRegWriteData[22]~3_combout\ <= NOT \Comb:vRegWriteData[22]~3_combout\;
\ALT_INV_Comb:vRegWriteData[22]~2_combout\ <= NOT \Comb:vRegWriteData[22]~2_combout\;
\ALT_INV_Comb:vRegWriteData[22]~1_combout\ <= NOT \Comb:vRegWriteData[22]~1_combout\;
\ALT_INV_Comb:vRegWriteData[20]~3_combout\ <= NOT \Comb:vRegWriteData[20]~3_combout\;
\ALT_INV_Comb:vRegWriteData[20]~2_combout\ <= NOT \Comb:vRegWriteData[20]~2_combout\;
\ALT_INV_Comb:vRegWriteData[20]~1_combout\ <= NOT \Comb:vRegWriteData[20]~1_combout\;
\ALT_INV_Comb:vRegWriteData[27]~3_combout\ <= NOT \Comb:vRegWriteData[27]~3_combout\;
\ALT_INV_Comb:vRegWriteData[27]~2_combout\ <= NOT \Comb:vRegWriteData[27]~2_combout\;
\ALT_INV_Comb:vRegWriteData[27]~1_combout\ <= NOT \Comb:vRegWriteData[27]~1_combout\;
\ALT_INV_Comb:vRegWriteData[25]~3_combout\ <= NOT \Comb:vRegWriteData[25]~3_combout\;
\ALT_INV_Comb:vRegWriteData[25]~2_combout\ <= NOT \Comb:vRegWriteData[25]~2_combout\;
\ALT_INV_Comb:vRegWriteData[25]~1_combout\ <= NOT \Comb:vRegWriteData[25]~1_combout\;
\ALT_INV_Comb:vRegWriteData[24]~4_combout\ <= NOT \Comb:vRegWriteData[24]~4_combout\;
\ALT_INV_Comb:vRegWriteData[24]~3_combout\ <= NOT \Comb:vRegWriteData[24]~3_combout\;
\ALT_INV_Comb:vRegWriteData[24]~2_combout\ <= NOT \Comb:vRegWriteData[24]~2_combout\;
\ALT_INV_Equal3~13_combout\ <= NOT \Equal3~13_combout\;
\ALT_INV_Equal3~11_combout\ <= NOT \Equal3~11_combout\;
\ALT_INV_Equal3~10_combout\ <= NOT \Equal3~10_combout\;
\ALT_INV_Selector23~7_combout\ <= NOT \Selector23~7_combout\;
\ALT_INV_Comb:vRegWriteData[31]~2_combout\ <= NOT \Comb:vRegWriteData[31]~2_combout\;
\ALT_INV_Comb:vRegWriteData[31]~1_combout\ <= NOT \Comb:vRegWriteData[31]~1_combout\;
\ALT_INV_Comb:vRegWriteData[30]~2_combout\ <= NOT \Comb:vRegWriteData[30]~2_combout\;
\ALT_INV_Comb:vRegWriteData[30]~1_combout\ <= NOT \Comb:vRegWriteData[30]~1_combout\;
\ALT_INV_Comb:vRegWriteData[29]~2_combout\ <= NOT \Comb:vRegWriteData[29]~2_combout\;
\ALT_INV_Comb:vRegWriteData[29]~1_combout\ <= NOT \Comb:vRegWriteData[29]~1_combout\;
\ALT_INV_Comb:vRegWriteData[28]~2_combout\ <= NOT \Comb:vRegWriteData[28]~2_combout\;
\ALT_INV_Comb:vRegWriteData[28]~1_combout\ <= NOT \Comb:vRegWriteData[28]~1_combout\;
\ALT_INV_Comb:vRegWriteData[26]~2_combout\ <= NOT \Comb:vRegWriteData[26]~2_combout\;
\ALT_INV_Comb:vRegWriteData[26]~1_combout\ <= NOT \Comb:vRegWriteData[26]~1_combout\;
\ALT_INV_vAluRes~35_combout\ <= NOT \vAluRes~35_combout\;
\ALT_INV_vAluRes~34_combout\ <= NOT \vAluRes~34_combout\;
\ALT_INV_vAluRes~33_combout\ <= NOT \vAluRes~33_combout\;
\ALT_INV_vAluRes~32_combout\ <= NOT \vAluRes~32_combout\;
\ALT_INV_vAluRes~31_combout\ <= NOT \vAluRes~31_combout\;
\ALT_INV_Equal3~9_combout\ <= NOT \Equal3~9_combout\;
\ALT_INV_Selector13~5_combout\ <= NOT \Selector13~5_combout\;
\ALT_INV_Selector13~4_combout\ <= NOT \Selector13~4_combout\;
\ALT_INV_Mux31~0_combout\ <= NOT \Mux31~0_combout\;
\ALT_INV_Selector0~0_combout\ <= NOT \Selector0~0_combout\;
\ALT_INV_ShiftLeft0~58_combout\ <= NOT \ShiftLeft0~58_combout\;
\ALT_INV_ShiftLeft0~57_combout\ <= NOT \ShiftLeft0~57_combout\;
\ALT_INV_Equal3~8_combout\ <= NOT \Equal3~8_combout\;
\ALT_INV_Equal3~6_combout\ <= NOT \Equal3~6_combout\;
\ALT_INV_Equal3~2_combout\ <= NOT \Equal3~2_combout\;
\ALT_INV_RegFile[26][23]~q\ <= NOT \RegFile[26][23]~q\;
\ALT_INV_RegFile[24][23]~q\ <= NOT \RegFile[24][23]~q\;
\ALT_INV_RegFile[27][23]~q\ <= NOT \RegFile[27][23]~q\;
\ALT_INV_RegFile[25][23]~q\ <= NOT \RegFile[25][23]~q\;
\ALT_INV_RegFile[18][23]~q\ <= NOT \RegFile[18][23]~q\;
\ALT_INV_RegFile[16][23]~q\ <= NOT \RegFile[16][23]~q\;
\ALT_INV_RegFile[19][23]~q\ <= NOT \RegFile[19][23]~q\;
\ALT_INV_RegFile[17][23]~q\ <= NOT \RegFile[17][23]~q\;
\ALT_INV_RegFile[10][23]~q\ <= NOT \RegFile[10][23]~q\;
\ALT_INV_RegFile[8][23]~q\ <= NOT \RegFile[8][23]~q\;
\ALT_INV_RegFile[11][23]~q\ <= NOT \RegFile[11][23]~q\;
\ALT_INV_RegFile[9][23]~q\ <= NOT \RegFile[9][23]~q\;
\ALT_INV_RegFile[26][22]~q\ <= NOT \RegFile[26][22]~q\;
\ALT_INV_RegFile[24][22]~q\ <= NOT \RegFile[24][22]~q\;
\ALT_INV_RegFile[27][22]~q\ <= NOT \RegFile[27][22]~q\;
\ALT_INV_RegFile[25][22]~q\ <= NOT \RegFile[25][22]~q\;
\ALT_INV_RegFile[18][22]~q\ <= NOT \RegFile[18][22]~q\;
\ALT_INV_RegFile[16][22]~q\ <= NOT \RegFile[16][22]~q\;
\ALT_INV_RegFile[19][22]~q\ <= NOT \RegFile[19][22]~q\;
\ALT_INV_RegFile[17][22]~q\ <= NOT \RegFile[17][22]~q\;
\ALT_INV_RegFile[10][22]~q\ <= NOT \RegFile[10][22]~q\;
\ALT_INV_RegFile[8][22]~q\ <= NOT \RegFile[8][22]~q\;
\ALT_INV_RegFile[11][22]~q\ <= NOT \RegFile[11][22]~q\;
\ALT_INV_RegFile[9][22]~q\ <= NOT \RegFile[9][22]~q\;
\ALT_INV_RegFile[26][21]~q\ <= NOT \RegFile[26][21]~q\;
\ALT_INV_RegFile[24][21]~q\ <= NOT \RegFile[24][21]~q\;
\ALT_INV_RegFile[27][21]~q\ <= NOT \RegFile[27][21]~q\;
\ALT_INV_RegFile[25][21]~q\ <= NOT \RegFile[25][21]~q\;
\ALT_INV_RegFile[18][21]~q\ <= NOT \RegFile[18][21]~q\;
\ALT_INV_RegFile[16][21]~q\ <= NOT \RegFile[16][21]~q\;
\ALT_INV_RegFile[19][21]~q\ <= NOT \RegFile[19][21]~q\;
\ALT_INV_RegFile[17][21]~q\ <= NOT \RegFile[17][21]~q\;
\ALT_INV_RegFile[10][21]~q\ <= NOT \RegFile[10][21]~q\;
\ALT_INV_RegFile[8][21]~q\ <= NOT \RegFile[8][21]~q\;
\ALT_INV_RegFile[11][21]~q\ <= NOT \RegFile[11][21]~q\;
\ALT_INV_RegFile[9][21]~q\ <= NOT \RegFile[9][21]~q\;
\ALT_INV_RegFile[26][20]~q\ <= NOT \RegFile[26][20]~q\;
\ALT_INV_RegFile[24][20]~q\ <= NOT \RegFile[24][20]~q\;
\ALT_INV_RegFile[27][20]~q\ <= NOT \RegFile[27][20]~q\;
\ALT_INV_RegFile[25][20]~q\ <= NOT \RegFile[25][20]~q\;
\ALT_INV_RegFile[18][20]~q\ <= NOT \RegFile[18][20]~q\;
\ALT_INV_RegFile[16][20]~q\ <= NOT \RegFile[16][20]~q\;
\ALT_INV_RegFile[19][20]~q\ <= NOT \RegFile[19][20]~q\;
\ALT_INV_RegFile[17][20]~q\ <= NOT \RegFile[17][20]~q\;
\ALT_INV_RegFile[10][20]~q\ <= NOT \RegFile[10][20]~q\;
\ALT_INV_RegFile[8][20]~q\ <= NOT \RegFile[8][20]~q\;
\ALT_INV_RegFile[11][20]~q\ <= NOT \RegFile[11][20]~q\;
\ALT_INV_RegFile[9][20]~q\ <= NOT \RegFile[9][20]~q\;
\ALT_INV_RegFile[26][19]~q\ <= NOT \RegFile[26][19]~q\;
\ALT_INV_RegFile[24][19]~q\ <= NOT \RegFile[24][19]~q\;
\ALT_INV_RegFile[27][19]~q\ <= NOT \RegFile[27][19]~q\;
\ALT_INV_RegFile[25][19]~q\ <= NOT \RegFile[25][19]~q\;
\ALT_INV_RegFile[18][19]~q\ <= NOT \RegFile[18][19]~q\;
\ALT_INV_RegFile[16][19]~q\ <= NOT \RegFile[16][19]~q\;
\ALT_INV_RegFile[19][19]~q\ <= NOT \RegFile[19][19]~q\;
\ALT_INV_RegFile[17][19]~q\ <= NOT \RegFile[17][19]~q\;
\ALT_INV_RegFile[10][19]~q\ <= NOT \RegFile[10][19]~q\;
\ALT_INV_RegFile[8][19]~q\ <= NOT \RegFile[8][19]~q\;
\ALT_INV_RegFile[11][19]~q\ <= NOT \RegFile[11][19]~q\;
\ALT_INV_RegFile[9][19]~q\ <= NOT \RegFile[9][19]~q\;
\ALT_INV_Comb:vRegWriteData[19]~0_combout\ <= NOT \Comb:vRegWriteData[19]~0_combout\;
\ALT_INV_RegFile[26][18]~q\ <= NOT \RegFile[26][18]~q\;
\ALT_INV_RegFile[24][18]~q\ <= NOT \RegFile[24][18]~q\;
\ALT_INV_RegFile[27][18]~q\ <= NOT \RegFile[27][18]~q\;
\ALT_INV_RegFile[25][18]~q\ <= NOT \RegFile[25][18]~q\;
\ALT_INV_RegFile[18][18]~q\ <= NOT \RegFile[18][18]~q\;
\ALT_INV_RegFile[16][18]~q\ <= NOT \RegFile[16][18]~q\;
\ALT_INV_RegFile[19][18]~q\ <= NOT \RegFile[19][18]~q\;
\ALT_INV_RegFile[17][18]~q\ <= NOT \RegFile[17][18]~q\;
\ALT_INV_RegFile[10][18]~q\ <= NOT \RegFile[10][18]~q\;
\ALT_INV_RegFile[8][18]~q\ <= NOT \RegFile[8][18]~q\;
\ALT_INV_RegFile[11][18]~q\ <= NOT \RegFile[11][18]~q\;
\ALT_INV_RegFile[9][18]~q\ <= NOT \RegFile[9][18]~q\;
\ALT_INV_RegFile[26][17]~q\ <= NOT \RegFile[26][17]~q\;
\ALT_INV_RegFile[24][17]~q\ <= NOT \RegFile[24][17]~q\;
\ALT_INV_RegFile[27][17]~q\ <= NOT \RegFile[27][17]~q\;
\ALT_INV_RegFile[25][17]~q\ <= NOT \RegFile[25][17]~q\;
\ALT_INV_RegFile[18][17]~q\ <= NOT \RegFile[18][17]~q\;
\ALT_INV_RegFile[16][17]~q\ <= NOT \RegFile[16][17]~q\;
\ALT_INV_RegFile[19][17]~q\ <= NOT \RegFile[19][17]~q\;
\ALT_INV_RegFile[17][17]~q\ <= NOT \RegFile[17][17]~q\;
\ALT_INV_RegFile[10][17]~q\ <= NOT \RegFile[10][17]~q\;
\ALT_INV_RegFile[8][17]~q\ <= NOT \RegFile[8][17]~q\;
\ALT_INV_RegFile[11][17]~q\ <= NOT \RegFile[11][17]~q\;
\ALT_INV_RegFile[9][17]~q\ <= NOT \RegFile[9][17]~q\;
\ALT_INV_RegFile[26][16]~q\ <= NOT \RegFile[26][16]~q\;
\ALT_INV_RegFile[24][16]~q\ <= NOT \RegFile[24][16]~q\;
\ALT_INV_RegFile[27][16]~q\ <= NOT \RegFile[27][16]~q\;
\ALT_INV_RegFile[25][16]~q\ <= NOT \RegFile[25][16]~q\;
\ALT_INV_RegFile[18][16]~q\ <= NOT \RegFile[18][16]~q\;
\ALT_INV_RegFile[16][16]~q\ <= NOT \RegFile[16][16]~q\;
\ALT_INV_RegFile[19][16]~q\ <= NOT \RegFile[19][16]~q\;
\ALT_INV_RegFile[17][16]~q\ <= NOT \RegFile[17][16]~q\;
\ALT_INV_RegFile[10][16]~q\ <= NOT \RegFile[10][16]~q\;
\ALT_INV_RegFile[8][16]~q\ <= NOT \RegFile[8][16]~q\;
\ALT_INV_RegFile[11][16]~q\ <= NOT \RegFile[11][16]~q\;
\ALT_INV_RegFile[9][16]~q\ <= NOT \RegFile[9][16]~q\;
\ALT_INV_Comb:vRegWriteData[24]~1_combout\ <= NOT \Comb:vRegWriteData[24]~1_combout\;
\ALT_INV_RegFile[26][7]~q\ <= NOT \RegFile[26][7]~q\;
\ALT_INV_RegFile[24][7]~q\ <= NOT \RegFile[24][7]~q\;
\ALT_INV_RegFile[27][7]~q\ <= NOT \RegFile[27][7]~q\;
\ALT_INV_RegFile[25][7]~q\ <= NOT \RegFile[25][7]~q\;
\ALT_INV_RegFile[18][7]~q\ <= NOT \RegFile[18][7]~q\;
\ALT_INV_RegFile[16][7]~q\ <= NOT \RegFile[16][7]~q\;
\ALT_INV_RegFile[19][7]~q\ <= NOT \RegFile[19][7]~q\;
\ALT_INV_RegFile[17][7]~q\ <= NOT \RegFile[17][7]~q\;
\ALT_INV_RegFile[10][7]~q\ <= NOT \RegFile[10][7]~q\;
\ALT_INV_RegFile[8][7]~q\ <= NOT \RegFile[8][7]~q\;
\ALT_INV_RegFile[11][7]~q\ <= NOT \RegFile[11][7]~q\;
\ALT_INV_RegFile[9][7]~q\ <= NOT \RegFile[9][7]~q\;
\ALT_INV_RegFile[26][15]~q\ <= NOT \RegFile[26][15]~q\;
\ALT_INV_RegFile[24][15]~q\ <= NOT \RegFile[24][15]~q\;
\ALT_INV_RegFile[27][15]~q\ <= NOT \RegFile[27][15]~q\;
\ALT_INV_RegFile[25][15]~q\ <= NOT \RegFile[25][15]~q\;
\ALT_INV_RegFile[18][15]~q\ <= NOT \RegFile[18][15]~q\;
\ALT_INV_RegFile[16][15]~q\ <= NOT \RegFile[16][15]~q\;
\ALT_INV_RegFile[19][15]~q\ <= NOT \RegFile[19][15]~q\;
\ALT_INV_RegFile[17][15]~q\ <= NOT \RegFile[17][15]~q\;
\ALT_INV_RegFile[10][15]~q\ <= NOT \RegFile[10][15]~q\;
\ALT_INV_RegFile[8][15]~q\ <= NOT \RegFile[8][15]~q\;
\ALT_INV_RegFile[11][15]~q\ <= NOT \RegFile[11][15]~q\;
\ALT_INV_RegFile[9][15]~q\ <= NOT \RegFile[9][15]~q\;
\ALT_INV_RegFile[26][31]~q\ <= NOT \RegFile[26][31]~q\;
\ALT_INV_RegFile[24][31]~q\ <= NOT \RegFile[24][31]~q\;
\ALT_INV_RegFile[27][31]~q\ <= NOT \RegFile[27][31]~q\;
\ALT_INV_RegFile[25][31]~q\ <= NOT \RegFile[25][31]~q\;
\ALT_INV_RegFile[18][31]~q\ <= NOT \RegFile[18][31]~q\;
\ALT_INV_RegFile[16][31]~q\ <= NOT \RegFile[16][31]~q\;
\ALT_INV_RegFile[19][31]~q\ <= NOT \RegFile[19][31]~q\;
\ALT_INV_RegFile[17][31]~q\ <= NOT \RegFile[17][31]~q\;
\ALT_INV_RegFile[10][31]~q\ <= NOT \RegFile[10][31]~q\;
\ALT_INV_RegFile[8][31]~q\ <= NOT \RegFile[8][31]~q\;
\ALT_INV_RegFile[11][31]~q\ <= NOT \RegFile[11][31]~q\;
\ALT_INV_RegFile[9][31]~q\ <= NOT \RegFile[9][31]~q\;
\ALT_INV_RegFile[26][6]~q\ <= NOT \RegFile[26][6]~q\;
\ALT_INV_RegFile[24][6]~q\ <= NOT \RegFile[24][6]~q\;
\ALT_INV_RegFile[27][6]~q\ <= NOT \RegFile[27][6]~q\;
\ALT_INV_RegFile[25][6]~q\ <= NOT \RegFile[25][6]~q\;
\ALT_INV_RegFile[18][6]~q\ <= NOT \RegFile[18][6]~q\;
\ALT_INV_RegFile[16][6]~q\ <= NOT \RegFile[16][6]~q\;
\ALT_INV_RegFile[19][6]~q\ <= NOT \RegFile[19][6]~q\;
\ALT_INV_RegFile[17][6]~q\ <= NOT \RegFile[17][6]~q\;
\ALT_INV_RegFile[10][6]~q\ <= NOT \RegFile[10][6]~q\;
\ALT_INV_RegFile[8][6]~q\ <= NOT \RegFile[8][6]~q\;
\ALT_INV_RegFile[11][6]~q\ <= NOT \RegFile[11][6]~q\;
\ALT_INV_RegFile[9][6]~q\ <= NOT \RegFile[9][6]~q\;
\ALT_INV_RegFile[26][14]~q\ <= NOT \RegFile[26][14]~q\;
\ALT_INV_RegFile[24][14]~q\ <= NOT \RegFile[24][14]~q\;
\ALT_INV_RegFile[27][14]~q\ <= NOT \RegFile[27][14]~q\;
\ALT_INV_RegFile[25][14]~q\ <= NOT \RegFile[25][14]~q\;
\ALT_INV_RegFile[18][14]~q\ <= NOT \RegFile[18][14]~q\;
\ALT_INV_RegFile[16][14]~q\ <= NOT \RegFile[16][14]~q\;
\ALT_INV_RegFile[19][14]~q\ <= NOT \RegFile[19][14]~q\;
\ALT_INV_RegFile[17][14]~q\ <= NOT \RegFile[17][14]~q\;
\ALT_INV_RegFile[10][14]~q\ <= NOT \RegFile[10][14]~q\;
\ALT_INV_RegFile[8][14]~q\ <= NOT \RegFile[8][14]~q\;
\ALT_INV_RegFile[11][14]~q\ <= NOT \RegFile[11][14]~q\;
\ALT_INV_RegFile[9][14]~q\ <= NOT \RegFile[9][14]~q\;
\ALT_INV_RegFile[26][30]~q\ <= NOT \RegFile[26][30]~q\;
\ALT_INV_RegFile[24][30]~q\ <= NOT \RegFile[24][30]~q\;
\ALT_INV_RegFile[27][30]~q\ <= NOT \RegFile[27][30]~q\;
\ALT_INV_RegFile[25][30]~q\ <= NOT \RegFile[25][30]~q\;
\ALT_INV_RegFile[18][30]~q\ <= NOT \RegFile[18][30]~q\;
\ALT_INV_RegFile[16][30]~q\ <= NOT \RegFile[16][30]~q\;
\ALT_INV_RegFile[19][30]~q\ <= NOT \RegFile[19][30]~q\;
\ALT_INV_RegFile[17][30]~q\ <= NOT \RegFile[17][30]~q\;
\ALT_INV_RegFile[10][30]~q\ <= NOT \RegFile[10][30]~q\;
\ALT_INV_RegFile[8][30]~q\ <= NOT \RegFile[8][30]~q\;
\ALT_INV_RegFile[11][30]~q\ <= NOT \RegFile[11][30]~q\;
\ALT_INV_RegFile[9][30]~q\ <= NOT \RegFile[9][30]~q\;
\ALT_INV_RegFile[26][5]~q\ <= NOT \RegFile[26][5]~q\;
\ALT_INV_RegFile[24][5]~q\ <= NOT \RegFile[24][5]~q\;
\ALT_INV_RegFile[27][5]~q\ <= NOT \RegFile[27][5]~q\;
\ALT_INV_RegFile[25][5]~q\ <= NOT \RegFile[25][5]~q\;
\ALT_INV_RegFile[18][5]~q\ <= NOT \RegFile[18][5]~q\;
\ALT_INV_RegFile[16][5]~q\ <= NOT \RegFile[16][5]~q\;
\ALT_INV_RegFile[19][5]~q\ <= NOT \RegFile[19][5]~q\;
\ALT_INV_RegFile[17][5]~q\ <= NOT \RegFile[17][5]~q\;
\ALT_INV_RegFile[10][5]~q\ <= NOT \RegFile[10][5]~q\;
\ALT_INV_RegFile[8][5]~q\ <= NOT \RegFile[8][5]~q\;
\ALT_INV_RegFile[11][5]~q\ <= NOT \RegFile[11][5]~q\;
\ALT_INV_RegFile[9][5]~q\ <= NOT \RegFile[9][5]~q\;
\ALT_INV_RegFile[26][13]~q\ <= NOT \RegFile[26][13]~q\;
\ALT_INV_RegFile[24][13]~q\ <= NOT \RegFile[24][13]~q\;
\ALT_INV_RegFile[27][13]~q\ <= NOT \RegFile[27][13]~q\;
\ALT_INV_RegFile[25][13]~q\ <= NOT \RegFile[25][13]~q\;
\ALT_INV_RegFile[18][13]~q\ <= NOT \RegFile[18][13]~q\;
\ALT_INV_RegFile[16][13]~q\ <= NOT \RegFile[16][13]~q\;
\ALT_INV_RegFile[19][13]~q\ <= NOT \RegFile[19][13]~q\;
\ALT_INV_RegFile[17][13]~q\ <= NOT \RegFile[17][13]~q\;
\ALT_INV_RegFile[10][13]~q\ <= NOT \RegFile[10][13]~q\;
\ALT_INV_RegFile[8][13]~q\ <= NOT \RegFile[8][13]~q\;
\ALT_INV_RegFile[11][13]~q\ <= NOT \RegFile[11][13]~q\;
\ALT_INV_RegFile[9][13]~q\ <= NOT \RegFile[9][13]~q\;
\ALT_INV_RegFile[26][29]~q\ <= NOT \RegFile[26][29]~q\;
\ALT_INV_RegFile[24][29]~q\ <= NOT \RegFile[24][29]~q\;
\ALT_INV_RegFile[27][29]~q\ <= NOT \RegFile[27][29]~q\;
\ALT_INV_RegFile[25][29]~q\ <= NOT \RegFile[25][29]~q\;
\ALT_INV_RegFile[18][29]~q\ <= NOT \RegFile[18][29]~q\;
\ALT_INV_RegFile[16][29]~q\ <= NOT \RegFile[16][29]~q\;
\ALT_INV_RegFile[19][29]~q\ <= NOT \RegFile[19][29]~q\;
\ALT_INV_RegFile[17][29]~q\ <= NOT \RegFile[17][29]~q\;
\ALT_INV_RegFile[10][29]~q\ <= NOT \RegFile[10][29]~q\;
\ALT_INV_RegFile[8][29]~q\ <= NOT \RegFile[8][29]~q\;
\ALT_INV_RegFile[11][29]~q\ <= NOT \RegFile[11][29]~q\;
\ALT_INV_RegFile[9][29]~q\ <= NOT \RegFile[9][29]~q\;
\ALT_INV_RegFile[26][4]~q\ <= NOT \RegFile[26][4]~q\;
\ALT_INV_RegFile[24][4]~q\ <= NOT \RegFile[24][4]~q\;
\ALT_INV_RegFile[27][4]~q\ <= NOT \RegFile[27][4]~q\;
\ALT_INV_RegFile[25][4]~q\ <= NOT \RegFile[25][4]~q\;
\ALT_INV_RegFile[18][4]~q\ <= NOT \RegFile[18][4]~q\;
\ALT_INV_RegFile[16][4]~q\ <= NOT \RegFile[16][4]~q\;
\ALT_INV_RegFile[19][4]~q\ <= NOT \RegFile[19][4]~q\;
\ALT_INV_RegFile[17][4]~q\ <= NOT \RegFile[17][4]~q\;
\ALT_INV_RegFile[10][4]~q\ <= NOT \RegFile[10][4]~q\;
\ALT_INV_RegFile[8][4]~q\ <= NOT \RegFile[8][4]~q\;
\ALT_INV_RegFile[11][4]~q\ <= NOT \RegFile[11][4]~q\;
\ALT_INV_RegFile[9][4]~q\ <= NOT \RegFile[9][4]~q\;
\ALT_INV_RegFile[26][12]~q\ <= NOT \RegFile[26][12]~q\;
\ALT_INV_RegFile[24][12]~q\ <= NOT \RegFile[24][12]~q\;
\ALT_INV_RegFile[27][12]~q\ <= NOT \RegFile[27][12]~q\;
\ALT_INV_RegFile[25][12]~q\ <= NOT \RegFile[25][12]~q\;
\ALT_INV_RegFile[18][12]~q\ <= NOT \RegFile[18][12]~q\;
\ALT_INV_RegFile[16][12]~q\ <= NOT \RegFile[16][12]~q\;
\ALT_INV_RegFile[19][12]~q\ <= NOT \RegFile[19][12]~q\;
\ALT_INV_RegFile[17][12]~q\ <= NOT \RegFile[17][12]~q\;
\ALT_INV_RegFile[10][12]~q\ <= NOT \RegFile[10][12]~q\;
\ALT_INV_RegFile[8][12]~q\ <= NOT \RegFile[8][12]~q\;
\ALT_INV_RegFile[11][12]~q\ <= NOT \RegFile[11][12]~q\;
\ALT_INV_RegFile[9][12]~q\ <= NOT \RegFile[9][12]~q\;
\ALT_INV_RegFile[26][28]~q\ <= NOT \RegFile[26][28]~q\;
\ALT_INV_RegFile[24][28]~q\ <= NOT \RegFile[24][28]~q\;
\ALT_INV_RegFile[27][28]~q\ <= NOT \RegFile[27][28]~q\;
\ALT_INV_RegFile[25][28]~q\ <= NOT \RegFile[25][28]~q\;
\ALT_INV_RegFile[18][28]~q\ <= NOT \RegFile[18][28]~q\;
\ALT_INV_RegFile[16][28]~q\ <= NOT \RegFile[16][28]~q\;
\ALT_INV_RegFile[19][28]~q\ <= NOT \RegFile[19][28]~q\;
\ALT_INV_RegFile[17][28]~q\ <= NOT \RegFile[17][28]~q\;
\ALT_INV_RegFile[10][28]~q\ <= NOT \RegFile[10][28]~q\;
\ALT_INV_RegFile[8][28]~q\ <= NOT \RegFile[8][28]~q\;
\ALT_INV_RegFile[11][28]~q\ <= NOT \RegFile[11][28]~q\;
\ALT_INV_RegFile[9][28]~q\ <= NOT \RegFile[9][28]~q\;
\ALT_INV_RegFile[26][3]~q\ <= NOT \RegFile[26][3]~q\;
\ALT_INV_RegFile[24][3]~q\ <= NOT \RegFile[24][3]~q\;
\ALT_INV_RegFile[27][3]~q\ <= NOT \RegFile[27][3]~q\;
\ALT_INV_RegFile[25][3]~q\ <= NOT \RegFile[25][3]~q\;
\ALT_INV_RegFile[18][3]~q\ <= NOT \RegFile[18][3]~q\;
\ALT_INV_RegFile[16][3]~q\ <= NOT \RegFile[16][3]~q\;
\ALT_INV_RegFile[19][3]~q\ <= NOT \RegFile[19][3]~q\;
\ALT_INV_RegFile[17][3]~q\ <= NOT \RegFile[17][3]~q\;
\ALT_INV_RegFile[10][3]~q\ <= NOT \RegFile[10][3]~q\;
\ALT_INV_RegFile[8][3]~q\ <= NOT \RegFile[8][3]~q\;
\ALT_INV_RegFile[11][3]~q\ <= NOT \RegFile[11][3]~q\;
\ALT_INV_RegFile[9][3]~q\ <= NOT \RegFile[9][3]~q\;
\ALT_INV_RegFile[26][11]~q\ <= NOT \RegFile[26][11]~q\;
\ALT_INV_RegFile[24][11]~q\ <= NOT \RegFile[24][11]~q\;
\ALT_INV_RegFile[27][11]~q\ <= NOT \RegFile[27][11]~q\;
\ALT_INV_RegFile[25][11]~q\ <= NOT \RegFile[25][11]~q\;
\ALT_INV_RegFile[18][11]~q\ <= NOT \RegFile[18][11]~q\;
\ALT_INV_RegFile[16][11]~q\ <= NOT \RegFile[16][11]~q\;
\ALT_INV_RegFile[19][11]~q\ <= NOT \RegFile[19][11]~q\;
\ALT_INV_RegFile[17][11]~q\ <= NOT \RegFile[17][11]~q\;
\ALT_INV_RegFile[10][11]~q\ <= NOT \RegFile[10][11]~q\;
\ALT_INV_RegFile[8][11]~q\ <= NOT \RegFile[8][11]~q\;
\ALT_INV_RegFile[11][11]~q\ <= NOT \RegFile[11][11]~q\;
\ALT_INV_RegFile[9][11]~q\ <= NOT \RegFile[9][11]~q\;
\ALT_INV_RegFile[26][27]~q\ <= NOT \RegFile[26][27]~q\;
\ALT_INV_RegFile[24][27]~q\ <= NOT \RegFile[24][27]~q\;
\ALT_INV_RegFile[27][27]~q\ <= NOT \RegFile[27][27]~q\;
\ALT_INV_RegFile[25][27]~q\ <= NOT \RegFile[25][27]~q\;
\ALT_INV_RegFile[18][27]~q\ <= NOT \RegFile[18][27]~q\;
\ALT_INV_RegFile[16][27]~q\ <= NOT \RegFile[16][27]~q\;
\ALT_INV_RegFile[19][27]~q\ <= NOT \RegFile[19][27]~q\;
\ALT_INV_RegFile[17][27]~q\ <= NOT \RegFile[17][27]~q\;
\ALT_INV_RegFile[10][27]~q\ <= NOT \RegFile[10][27]~q\;
\ALT_INV_RegFile[8][27]~q\ <= NOT \RegFile[8][27]~q\;
\ALT_INV_RegFile[11][27]~q\ <= NOT \RegFile[11][27]~q\;
\ALT_INV_RegFile[9][27]~q\ <= NOT \RegFile[9][27]~q\;
\ALT_INV_RegFile[26][2]~q\ <= NOT \RegFile[26][2]~q\;
\ALT_INV_RegFile[24][2]~q\ <= NOT \RegFile[24][2]~q\;
\ALT_INV_RegFile[27][2]~q\ <= NOT \RegFile[27][2]~q\;
\ALT_INV_RegFile[25][2]~q\ <= NOT \RegFile[25][2]~q\;
\ALT_INV_RegFile[18][2]~q\ <= NOT \RegFile[18][2]~q\;
\ALT_INV_RegFile[16][2]~q\ <= NOT \RegFile[16][2]~q\;
\ALT_INV_RegFile[19][2]~q\ <= NOT \RegFile[19][2]~q\;
\ALT_INV_RegFile[17][2]~q\ <= NOT \RegFile[17][2]~q\;
\ALT_INV_RegFile[10][2]~q\ <= NOT \RegFile[10][2]~q\;
\ALT_INV_RegFile[8][2]~q\ <= NOT \RegFile[8][2]~q\;
\ALT_INV_RegFile[11][2]~q\ <= NOT \RegFile[11][2]~q\;
\ALT_INV_RegFile[9][2]~q\ <= NOT \RegFile[9][2]~q\;
\ALT_INV_RegFile[26][10]~q\ <= NOT \RegFile[26][10]~q\;
\ALT_INV_RegFile[24][10]~q\ <= NOT \RegFile[24][10]~q\;
\ALT_INV_RegFile[27][10]~q\ <= NOT \RegFile[27][10]~q\;
\ALT_INV_RegFile[25][10]~q\ <= NOT \RegFile[25][10]~q\;
\ALT_INV_RegFile[18][10]~q\ <= NOT \RegFile[18][10]~q\;
\ALT_INV_RegFile[16][10]~q\ <= NOT \RegFile[16][10]~q\;
\ALT_INV_RegFile[19][10]~q\ <= NOT \RegFile[19][10]~q\;
\ALT_INV_RegFile[17][10]~q\ <= NOT \RegFile[17][10]~q\;
\ALT_INV_RegFile[10][10]~q\ <= NOT \RegFile[10][10]~q\;
\ALT_INV_RegFile[8][10]~q\ <= NOT \RegFile[8][10]~q\;
\ALT_INV_RegFile[11][10]~q\ <= NOT \RegFile[11][10]~q\;
\ALT_INV_RegFile[9][10]~q\ <= NOT \RegFile[9][10]~q\;
\ALT_INV_Comb:vRegWriteData[10]~0_combout\ <= NOT \Comb:vRegWriteData[10]~0_combout\;
\ALT_INV_RegFile[26][26]~q\ <= NOT \RegFile[26][26]~q\;
\ALT_INV_RegFile[24][26]~q\ <= NOT \RegFile[24][26]~q\;
\ALT_INV_RegFile[27][26]~q\ <= NOT \RegFile[27][26]~q\;
\ALT_INV_RegFile[25][26]~q\ <= NOT \RegFile[25][26]~q\;
\ALT_INV_RegFile[18][26]~q\ <= NOT \RegFile[18][26]~q\;
\ALT_INV_RegFile[16][26]~q\ <= NOT \RegFile[16][26]~q\;
\ALT_INV_RegFile[19][26]~q\ <= NOT \RegFile[19][26]~q\;
\ALT_INV_RegFile[17][26]~q\ <= NOT \RegFile[17][26]~q\;
\ALT_INV_RegFile[10][26]~q\ <= NOT \RegFile[10][26]~q\;
\ALT_INV_RegFile[8][26]~q\ <= NOT \RegFile[8][26]~q\;
\ALT_INV_RegFile[11][26]~q\ <= NOT \RegFile[11][26]~q\;
\ALT_INV_RegFile[9][26]~q\ <= NOT \RegFile[9][26]~q\;
\ALT_INV_RegFile[26][1]~q\ <= NOT \RegFile[26][1]~q\;
\ALT_INV_RegFile[24][1]~q\ <= NOT \RegFile[24][1]~q\;
\ALT_INV_RegFile[27][1]~q\ <= NOT \RegFile[27][1]~q\;
\ALT_INV_RegFile[25][1]~q\ <= NOT \RegFile[25][1]~q\;
\ALT_INV_RegFile[18][1]~q\ <= NOT \RegFile[18][1]~q\;
\ALT_INV_RegFile[16][1]~q\ <= NOT \RegFile[16][1]~q\;
\ALT_INV_RegFile[19][1]~q\ <= NOT \RegFile[19][1]~q\;
\ALT_INV_RegFile[17][1]~q\ <= NOT \RegFile[17][1]~q\;
\ALT_INV_RegFile[10][1]~q\ <= NOT \RegFile[10][1]~q\;
\ALT_INV_RegFile[8][1]~q\ <= NOT \RegFile[8][1]~q\;
\ALT_INV_RegFile[11][1]~q\ <= NOT \RegFile[11][1]~q\;
\ALT_INV_RegFile[9][1]~q\ <= NOT \RegFile[9][1]~q\;
\ALT_INV_RegFile[26][9]~q\ <= NOT \RegFile[26][9]~q\;
\ALT_INV_RegFile[24][9]~q\ <= NOT \RegFile[24][9]~q\;
\ALT_INV_RegFile[27][9]~q\ <= NOT \RegFile[27][9]~q\;
\ALT_INV_RegFile[25][9]~q\ <= NOT \RegFile[25][9]~q\;
\ALT_INV_RegFile[18][9]~q\ <= NOT \RegFile[18][9]~q\;
\ALT_INV_RegFile[16][9]~q\ <= NOT \RegFile[16][9]~q\;
\ALT_INV_RegFile[19][9]~q\ <= NOT \RegFile[19][9]~q\;
\ALT_INV_RegFile[17][9]~q\ <= NOT \RegFile[17][9]~q\;
\ALT_INV_RegFile[10][9]~q\ <= NOT \RegFile[10][9]~q\;
\ALT_INV_RegFile[8][9]~q\ <= NOT \RegFile[8][9]~q\;
\ALT_INV_RegFile[11][9]~q\ <= NOT \RegFile[11][9]~q\;
\ALT_INV_RegFile[9][9]~q\ <= NOT \RegFile[9][9]~q\;
\ALT_INV_RegFile[26][25]~q\ <= NOT \RegFile[26][25]~q\;
\ALT_INV_RegFile[24][25]~q\ <= NOT \RegFile[24][25]~q\;
\ALT_INV_RegFile[27][25]~q\ <= NOT \RegFile[27][25]~q\;
\ALT_INV_RegFile[25][25]~q\ <= NOT \RegFile[25][25]~q\;
\ALT_INV_RegFile[18][25]~q\ <= NOT \RegFile[18][25]~q\;
\ALT_INV_RegFile[16][25]~q\ <= NOT \RegFile[16][25]~q\;
\ALT_INV_RegFile[19][25]~q\ <= NOT \RegFile[19][25]~q\;
\ALT_INV_RegFile[17][25]~q\ <= NOT \RegFile[17][25]~q\;
\ALT_INV_RegFile[10][25]~q\ <= NOT \RegFile[10][25]~q\;
\ALT_INV_RegFile[8][25]~q\ <= NOT \RegFile[8][25]~q\;
\ALT_INV_RegFile[11][25]~q\ <= NOT \RegFile[11][25]~q\;
\ALT_INV_RegFile[9][25]~q\ <= NOT \RegFile[9][25]~q\;
\ALT_INV_RegFile[26][0]~q\ <= NOT \RegFile[26][0]~q\;
\ALT_INV_RegFile[24][0]~q\ <= NOT \RegFile[24][0]~q\;
\ALT_INV_RegFile[27][0]~q\ <= NOT \RegFile[27][0]~q\;
\ALT_INV_RegFile[25][0]~q\ <= NOT \RegFile[25][0]~q\;
\ALT_INV_RegFile[18][0]~q\ <= NOT \RegFile[18][0]~q\;
\ALT_INV_RegFile[16][0]~q\ <= NOT \RegFile[16][0]~q\;
\ALT_INV_RegFile[19][0]~q\ <= NOT \RegFile[19][0]~q\;
\ALT_INV_RegFile[17][0]~q\ <= NOT \RegFile[17][0]~q\;
\ALT_INV_RegFile[10][0]~q\ <= NOT \RegFile[10][0]~q\;
\ALT_INV_RegFile[8][0]~q\ <= NOT \RegFile[8][0]~q\;
\ALT_INV_RegFile[11][0]~q\ <= NOT \RegFile[11][0]~q\;
\ALT_INV_RegFile[9][0]~q\ <= NOT \RegFile[9][0]~q\;
\ALT_INV_Comb:vRegWriteData[0]~0_combout\ <= NOT \Comb:vRegWriteData[0]~0_combout\;
\ALT_INV_RegFile[26][8]~q\ <= NOT \RegFile[26][8]~q\;
\ALT_INV_RegFile[24][8]~q\ <= NOT \RegFile[24][8]~q\;
\ALT_INV_RegFile[27][8]~q\ <= NOT \RegFile[27][8]~q\;
\ALT_INV_RegFile[25][8]~q\ <= NOT \RegFile[25][8]~q\;
\ALT_INV_RegFile[18][8]~q\ <= NOT \RegFile[18][8]~q\;
\ALT_INV_RegFile[16][8]~q\ <= NOT \RegFile[16][8]~q\;
\ALT_INV_RegFile[19][8]~q\ <= NOT \RegFile[19][8]~q\;
\ALT_INV_RegFile[17][8]~q\ <= NOT \RegFile[17][8]~q\;
\ALT_INV_RegFile[10][8]~q\ <= NOT \RegFile[10][8]~q\;
\ALT_INV_RegFile[8][8]~q\ <= NOT \RegFile[8][8]~q\;
\ALT_INV_RegFile[11][8]~q\ <= NOT \RegFile[11][8]~q\;
\ALT_INV_RegFile[9][8]~q\ <= NOT \RegFile[9][8]~q\;
\ALT_INV_RegFile[26][24]~q\ <= NOT \RegFile[26][24]~q\;
\ALT_INV_RegFile[24][24]~q\ <= NOT \RegFile[24][24]~q\;
\ALT_INV_RegFile[27][24]~q\ <= NOT \RegFile[27][24]~q\;
\ALT_INV_RegFile[25][24]~q\ <= NOT \RegFile[25][24]~q\;
\ALT_INV_RegFile[18][24]~q\ <= NOT \RegFile[18][24]~q\;
\ALT_INV_RegFile[16][24]~q\ <= NOT \RegFile[16][24]~q\;
\ALT_INV_RegFile[19][24]~q\ <= NOT \RegFile[19][24]~q\;
\ALT_INV_RegFile[17][24]~q\ <= NOT \RegFile[17][24]~q\;
\ALT_INV_RegFile[10][24]~q\ <= NOT \RegFile[10][24]~q\;
\ALT_INV_RegFile[8][24]~q\ <= NOT \RegFile[8][24]~q\;
\ALT_INV_RegFile[11][24]~q\ <= NOT \RegFile[11][24]~q\;
\ALT_INV_RegFile[9][24]~q\ <= NOT \RegFile[9][24]~q\;
\ALT_INV_R.regWriteEn~1_combout\ <= NOT \R.regWriteEn~1_combout\;
\ALT_INV_R.regWriteEn~0_combout\ <= NOT \R.regWriteEn~0_combout\;
\ALT_INV_NxR~15_combout\ <= NOT \NxR~15_combout\;
\ALT_INV_Mux50~0_combout\ <= NOT \Mux50~0_combout\;
\ALT_INV_Mux34~0_combout\ <= NOT \Mux34~0_combout\;
\ALT_INV_Mux11~0_combout\ <= NOT \Mux11~0_combout\;
\ALT_INV_NxR~10_combout\ <= NOT \NxR~10_combout\;
\ALT_INV_Mux44~0_combout\ <= NOT \Mux44~0_combout\;
\ALT_INV_NxR~9_combout\ <= NOT \NxR~9_combout\;
\ALT_INV_Mux58~0_combout\ <= NOT \Mux58~0_combout\;
\ALT_INV_R.statusReg\(2) <= NOT \R.statusReg\(2);
\ALT_INV_R.statusReg\(1) <= NOT \R.statusReg\(1);
\ALT_INV_R.ctrlState.CheckJump~q\ <= NOT \R.ctrlState.CheckJump~q\;
\ALT_INV_RegFile[30][23]~q\ <= NOT \RegFile[30][23]~q\;
\ALT_INV_RegFile[28][23]~q\ <= NOT \RegFile[28][23]~q\;
\ALT_INV_RegFile[31][23]~q\ <= NOT \RegFile[31][23]~q\;
\ALT_INV_RegFile[29][23]~q\ <= NOT \RegFile[29][23]~q\;
\ALT_INV_RegFile[22][23]~q\ <= NOT \RegFile[22][23]~q\;
\ALT_INV_RegFile[20][23]~q\ <= NOT \RegFile[20][23]~q\;
\ALT_INV_RegFile[23][23]~q\ <= NOT \RegFile[23][23]~q\;
\ALT_INV_RegFile[21][23]~q\ <= NOT \RegFile[21][23]~q\;
\ALT_INV_RegFile[14][23]~q\ <= NOT \RegFile[14][23]~q\;
\ALT_INV_RegFile[12][23]~q\ <= NOT \RegFile[12][23]~q\;
\ALT_INV_RegFile[15][23]~q\ <= NOT \RegFile[15][23]~q\;
\ALT_INV_RegFile[13][23]~q\ <= NOT \RegFile[13][23]~q\;
\ALT_INV_RegFile[30][22]~q\ <= NOT \RegFile[30][22]~q\;
\ALT_INV_RegFile[28][22]~q\ <= NOT \RegFile[28][22]~q\;
\ALT_INV_RegFile[31][22]~q\ <= NOT \RegFile[31][22]~q\;
\ALT_INV_RegFile[29][22]~q\ <= NOT \RegFile[29][22]~q\;
\ALT_INV_RegFile[22][22]~q\ <= NOT \RegFile[22][22]~q\;
\ALT_INV_RegFile[20][22]~q\ <= NOT \RegFile[20][22]~q\;
\ALT_INV_RegFile[23][22]~q\ <= NOT \RegFile[23][22]~q\;
\ALT_INV_RegFile[21][22]~q\ <= NOT \RegFile[21][22]~q\;
\ALT_INV_RegFile[14][22]~q\ <= NOT \RegFile[14][22]~q\;
\ALT_INV_RegFile[12][22]~q\ <= NOT \RegFile[12][22]~q\;
\ALT_INV_RegFile[15][22]~q\ <= NOT \RegFile[15][22]~q\;
\ALT_INV_RegFile[13][22]~q\ <= NOT \RegFile[13][22]~q\;
\ALT_INV_RegFile[30][21]~q\ <= NOT \RegFile[30][21]~q\;
\ALT_INV_RegFile[28][21]~q\ <= NOT \RegFile[28][21]~q\;
\ALT_INV_RegFile[31][21]~q\ <= NOT \RegFile[31][21]~q\;
\ALT_INV_RegFile[29][21]~q\ <= NOT \RegFile[29][21]~q\;
\ALT_INV_RegFile[22][21]~q\ <= NOT \RegFile[22][21]~q\;
\ALT_INV_RegFile[20][21]~q\ <= NOT \RegFile[20][21]~q\;
\ALT_INV_RegFile[23][21]~q\ <= NOT \RegFile[23][21]~q\;
\ALT_INV_RegFile[21][21]~q\ <= NOT \RegFile[21][21]~q\;
\ALT_INV_RegFile[14][21]~q\ <= NOT \RegFile[14][21]~q\;
\ALT_INV_RegFile[12][21]~q\ <= NOT \RegFile[12][21]~q\;
\ALT_INV_RegFile[15][21]~q\ <= NOT \RegFile[15][21]~q\;
\ALT_INV_RegFile[13][21]~q\ <= NOT \RegFile[13][21]~q\;
\ALT_INV_RegFile[30][20]~q\ <= NOT \RegFile[30][20]~q\;
\ALT_INV_RegFile[28][20]~q\ <= NOT \RegFile[28][20]~q\;
\ALT_INV_RegFile[31][20]~q\ <= NOT \RegFile[31][20]~q\;
\ALT_INV_RegFile[29][20]~q\ <= NOT \RegFile[29][20]~q\;
\ALT_INV_RegFile[22][20]~q\ <= NOT \RegFile[22][20]~q\;
\ALT_INV_RegFile[20][20]~q\ <= NOT \RegFile[20][20]~q\;
\ALT_INV_RegFile[23][20]~q\ <= NOT \RegFile[23][20]~q\;
\ALT_INV_RegFile[21][20]~q\ <= NOT \RegFile[21][20]~q\;
\ALT_INV_RegFile[14][20]~q\ <= NOT \RegFile[14][20]~q\;
\ALT_INV_RegFile[12][20]~q\ <= NOT \RegFile[12][20]~q\;
\ALT_INV_RegFile[15][20]~q\ <= NOT \RegFile[15][20]~q\;
\ALT_INV_RegFile[13][20]~q\ <= NOT \RegFile[13][20]~q\;
\ALT_INV_RegFile[30][19]~q\ <= NOT \RegFile[30][19]~q\;
\ALT_INV_RegFile[28][19]~q\ <= NOT \RegFile[28][19]~q\;
\ALT_INV_RegFile[31][19]~q\ <= NOT \RegFile[31][19]~q\;
\ALT_INV_RegFile[29][19]~q\ <= NOT \RegFile[29][19]~q\;
\ALT_INV_RegFile[22][19]~q\ <= NOT \RegFile[22][19]~q\;
\ALT_INV_RegFile[20][19]~q\ <= NOT \RegFile[20][19]~q\;
\ALT_INV_RegFile[23][19]~q\ <= NOT \RegFile[23][19]~q\;
\ALT_INV_RegFile[21][19]~q\ <= NOT \RegFile[21][19]~q\;
\ALT_INV_RegFile[14][19]~q\ <= NOT \RegFile[14][19]~q\;
\ALT_INV_RegFile[12][19]~q\ <= NOT \RegFile[12][19]~q\;
\ALT_INV_RegFile[15][19]~q\ <= NOT \RegFile[15][19]~q\;
\ALT_INV_RegFile[13][19]~q\ <= NOT \RegFile[13][19]~q\;
\ALT_INV_RegFile[30][18]~q\ <= NOT \RegFile[30][18]~q\;
\ALT_INV_RegFile[28][18]~q\ <= NOT \RegFile[28][18]~q\;
\ALT_INV_RegFile[31][18]~q\ <= NOT \RegFile[31][18]~q\;
\ALT_INV_RegFile[29][18]~q\ <= NOT \RegFile[29][18]~q\;
\ALT_INV_RegFile[22][18]~q\ <= NOT \RegFile[22][18]~q\;
\ALT_INV_RegFile[20][18]~q\ <= NOT \RegFile[20][18]~q\;
\ALT_INV_RegFile[23][18]~q\ <= NOT \RegFile[23][18]~q\;
\ALT_INV_RegFile[21][18]~q\ <= NOT \RegFile[21][18]~q\;
\ALT_INV_RegFile[14][18]~q\ <= NOT \RegFile[14][18]~q\;
\ALT_INV_RegFile[12][18]~q\ <= NOT \RegFile[12][18]~q\;
\ALT_INV_RegFile[15][18]~q\ <= NOT \RegFile[15][18]~q\;
\ALT_INV_RegFile[13][18]~q\ <= NOT \RegFile[13][18]~q\;
\ALT_INV_RegFile[30][17]~q\ <= NOT \RegFile[30][17]~q\;
\ALT_INV_RegFile[28][17]~q\ <= NOT \RegFile[28][17]~q\;
\ALT_INV_RegFile[31][17]~q\ <= NOT \RegFile[31][17]~q\;
\ALT_INV_RegFile[29][17]~q\ <= NOT \RegFile[29][17]~q\;
\ALT_INV_RegFile[22][17]~q\ <= NOT \RegFile[22][17]~q\;
\ALT_INV_RegFile[20][17]~q\ <= NOT \RegFile[20][17]~q\;
\ALT_INV_RegFile[23][17]~q\ <= NOT \RegFile[23][17]~q\;
\ALT_INV_RegFile[21][17]~q\ <= NOT \RegFile[21][17]~q\;
\ALT_INV_RegFile[14][17]~q\ <= NOT \RegFile[14][17]~q\;
\ALT_INV_RegFile[12][17]~q\ <= NOT \RegFile[12][17]~q\;
\ALT_INV_RegFile[15][17]~q\ <= NOT \RegFile[15][17]~q\;
\ALT_INV_RegFile[13][17]~q\ <= NOT \RegFile[13][17]~q\;
\ALT_INV_RegFile[30][16]~q\ <= NOT \RegFile[30][16]~q\;
\ALT_INV_RegFile[28][16]~q\ <= NOT \RegFile[28][16]~q\;
\ALT_INV_RegFile[31][16]~q\ <= NOT \RegFile[31][16]~q\;
\ALT_INV_RegFile[29][16]~q\ <= NOT \RegFile[29][16]~q\;
\ALT_INV_RegFile[22][16]~q\ <= NOT \RegFile[22][16]~q\;
\ALT_INV_RegFile[20][16]~q\ <= NOT \RegFile[20][16]~q\;
\ALT_INV_RegFile[23][16]~q\ <= NOT \RegFile[23][16]~q\;
\ALT_INV_RegFile[21][16]~q\ <= NOT \RegFile[21][16]~q\;
\ALT_INV_RegFile[14][16]~q\ <= NOT \RegFile[14][16]~q\;
\ALT_INV_RegFile[12][16]~q\ <= NOT \RegFile[12][16]~q\;
\ALT_INV_RegFile[15][16]~q\ <= NOT \RegFile[15][16]~q\;
\ALT_INV_RegFile[13][16]~q\ <= NOT \RegFile[13][16]~q\;
\ALT_INV_RegFile[30][7]~q\ <= NOT \RegFile[30][7]~q\;
\ALT_INV_RegFile[28][7]~q\ <= NOT \RegFile[28][7]~q\;
\ALT_INV_RegFile[31][7]~q\ <= NOT \RegFile[31][7]~q\;
\ALT_INV_RegFile[29][7]~q\ <= NOT \RegFile[29][7]~q\;
\ALT_INV_RegFile[22][7]~q\ <= NOT \RegFile[22][7]~q\;
\ALT_INV_RegFile[20][7]~q\ <= NOT \RegFile[20][7]~q\;
\ALT_INV_RegFile[23][7]~q\ <= NOT \RegFile[23][7]~q\;
\ALT_INV_RegFile[21][7]~q\ <= NOT \RegFile[21][7]~q\;
\ALT_INV_RegFile[14][7]~q\ <= NOT \RegFile[14][7]~q\;
\ALT_INV_RegFile[12][7]~q\ <= NOT \RegFile[12][7]~q\;
\ALT_INV_RegFile[15][7]~q\ <= NOT \RegFile[15][7]~q\;
\ALT_INV_RegFile[13][7]~q\ <= NOT \RegFile[13][7]~q\;
\ALT_INV_RegFile[30][15]~q\ <= NOT \RegFile[30][15]~q\;
\ALT_INV_RegFile[28][15]~q\ <= NOT \RegFile[28][15]~q\;
\ALT_INV_RegFile[31][15]~q\ <= NOT \RegFile[31][15]~q\;
\ALT_INV_RegFile[29][15]~q\ <= NOT \RegFile[29][15]~q\;
\ALT_INV_RegFile[22][15]~q\ <= NOT \RegFile[22][15]~q\;
\ALT_INV_RegFile[20][15]~q\ <= NOT \RegFile[20][15]~q\;
\ALT_INV_RegFile[23][15]~q\ <= NOT \RegFile[23][15]~q\;
\ALT_INV_RegFile[21][15]~q\ <= NOT \RegFile[21][15]~q\;
\ALT_INV_RegFile[14][15]~q\ <= NOT \RegFile[14][15]~q\;
\ALT_INV_RegFile[12][15]~q\ <= NOT \RegFile[12][15]~q\;
\ALT_INV_RegFile[15][15]~q\ <= NOT \RegFile[15][15]~q\;
\ALT_INV_RegFile[13][15]~q\ <= NOT \RegFile[13][15]~q\;
\ALT_INV_RegFile[30][31]~q\ <= NOT \RegFile[30][31]~q\;
\ALT_INV_RegFile[28][31]~q\ <= NOT \RegFile[28][31]~q\;
\ALT_INV_RegFile[31][31]~q\ <= NOT \RegFile[31][31]~q\;
\ALT_INV_RegFile[29][31]~q\ <= NOT \RegFile[29][31]~q\;
\ALT_INV_RegFile[22][31]~q\ <= NOT \RegFile[22][31]~q\;
\ALT_INV_RegFile[20][31]~q\ <= NOT \RegFile[20][31]~q\;
\ALT_INV_RegFile[23][31]~q\ <= NOT \RegFile[23][31]~q\;
\ALT_INV_RegFile[21][31]~q\ <= NOT \RegFile[21][31]~q\;
\ALT_INV_RegFile[14][31]~q\ <= NOT \RegFile[14][31]~q\;
\ALT_INV_RegFile[12][31]~q\ <= NOT \RegFile[12][31]~q\;
\ALT_INV_RegFile[15][31]~q\ <= NOT \RegFile[15][31]~q\;
\ALT_INV_RegFile[13][31]~q\ <= NOT \RegFile[13][31]~q\;
\ALT_INV_RegFile[30][6]~q\ <= NOT \RegFile[30][6]~q\;
\ALT_INV_RegFile[28][6]~q\ <= NOT \RegFile[28][6]~q\;
\ALT_INV_RegFile[31][6]~q\ <= NOT \RegFile[31][6]~q\;
\ALT_INV_RegFile[29][6]~q\ <= NOT \RegFile[29][6]~q\;
\ALT_INV_RegFile[22][6]~q\ <= NOT \RegFile[22][6]~q\;
\ALT_INV_RegFile[20][6]~q\ <= NOT \RegFile[20][6]~q\;
\ALT_INV_RegFile[23][6]~q\ <= NOT \RegFile[23][6]~q\;
\ALT_INV_RegFile[21][6]~q\ <= NOT \RegFile[21][6]~q\;
\ALT_INV_RegFile[14][6]~q\ <= NOT \RegFile[14][6]~q\;
\ALT_INV_RegFile[12][6]~q\ <= NOT \RegFile[12][6]~q\;
\ALT_INV_RegFile[15][6]~q\ <= NOT \RegFile[15][6]~q\;
\ALT_INV_RegFile[13][6]~q\ <= NOT \RegFile[13][6]~q\;
\ALT_INV_RegFile[30][14]~q\ <= NOT \RegFile[30][14]~q\;
\ALT_INV_RegFile[28][14]~q\ <= NOT \RegFile[28][14]~q\;
\ALT_INV_RegFile[31][14]~q\ <= NOT \RegFile[31][14]~q\;
\ALT_INV_RegFile[29][14]~q\ <= NOT \RegFile[29][14]~q\;
\ALT_INV_RegFile[22][14]~q\ <= NOT \RegFile[22][14]~q\;
\ALT_INV_RegFile[20][14]~q\ <= NOT \RegFile[20][14]~q\;
\ALT_INV_RegFile[23][14]~q\ <= NOT \RegFile[23][14]~q\;
\ALT_INV_RegFile[21][14]~q\ <= NOT \RegFile[21][14]~q\;
\ALT_INV_RegFile[14][14]~q\ <= NOT \RegFile[14][14]~q\;
\ALT_INV_RegFile[12][14]~q\ <= NOT \RegFile[12][14]~q\;
\ALT_INV_RegFile[15][14]~q\ <= NOT \RegFile[15][14]~q\;
\ALT_INV_RegFile[13][14]~q\ <= NOT \RegFile[13][14]~q\;
\ALT_INV_RegFile[30][30]~q\ <= NOT \RegFile[30][30]~q\;
\ALT_INV_RegFile[28][30]~q\ <= NOT \RegFile[28][30]~q\;
\ALT_INV_RegFile[31][30]~q\ <= NOT \RegFile[31][30]~q\;
\ALT_INV_RegFile[29][30]~q\ <= NOT \RegFile[29][30]~q\;
\ALT_INV_RegFile[22][30]~q\ <= NOT \RegFile[22][30]~q\;
\ALT_INV_RegFile[20][30]~q\ <= NOT \RegFile[20][30]~q\;
\ALT_INV_RegFile[23][30]~q\ <= NOT \RegFile[23][30]~q\;
\ALT_INV_RegFile[21][30]~q\ <= NOT \RegFile[21][30]~q\;
\ALT_INV_RegFile[14][30]~q\ <= NOT \RegFile[14][30]~q\;
\ALT_INV_RegFile[12][30]~q\ <= NOT \RegFile[12][30]~q\;
\ALT_INV_RegFile[15][30]~q\ <= NOT \RegFile[15][30]~q\;
\ALT_INV_RegFile[13][30]~q\ <= NOT \RegFile[13][30]~q\;
\ALT_INV_RegFile[30][5]~q\ <= NOT \RegFile[30][5]~q\;
\ALT_INV_RegFile[28][5]~q\ <= NOT \RegFile[28][5]~q\;
\ALT_INV_RegFile[31][5]~q\ <= NOT \RegFile[31][5]~q\;
\ALT_INV_RegFile[29][5]~q\ <= NOT \RegFile[29][5]~q\;
\ALT_INV_RegFile[22][5]~q\ <= NOT \RegFile[22][5]~q\;
\ALT_INV_RegFile[20][5]~q\ <= NOT \RegFile[20][5]~q\;
\ALT_INV_RegFile[23][5]~q\ <= NOT \RegFile[23][5]~q\;
\ALT_INV_RegFile[21][5]~q\ <= NOT \RegFile[21][5]~q\;
\ALT_INV_RegFile[14][5]~q\ <= NOT \RegFile[14][5]~q\;
\ALT_INV_RegFile[12][5]~q\ <= NOT \RegFile[12][5]~q\;
\ALT_INV_RegFile[15][5]~q\ <= NOT \RegFile[15][5]~q\;
\ALT_INV_RegFile[13][5]~q\ <= NOT \RegFile[13][5]~q\;
\ALT_INV_RegFile[30][13]~q\ <= NOT \RegFile[30][13]~q\;
\ALT_INV_RegFile[28][13]~q\ <= NOT \RegFile[28][13]~q\;
\ALT_INV_RegFile[31][13]~q\ <= NOT \RegFile[31][13]~q\;
\ALT_INV_RegFile[29][13]~q\ <= NOT \RegFile[29][13]~q\;
\ALT_INV_RegFile[22][13]~q\ <= NOT \RegFile[22][13]~q\;
\ALT_INV_RegFile[20][13]~q\ <= NOT \RegFile[20][13]~q\;
\ALT_INV_RegFile[23][13]~q\ <= NOT \RegFile[23][13]~q\;
\ALT_INV_RegFile[21][13]~q\ <= NOT \RegFile[21][13]~q\;
\ALT_INV_RegFile[14][13]~q\ <= NOT \RegFile[14][13]~q\;
\ALT_INV_RegFile[12][13]~q\ <= NOT \RegFile[12][13]~q\;
\ALT_INV_RegFile[15][13]~q\ <= NOT \RegFile[15][13]~q\;
\ALT_INV_RegFile[13][13]~q\ <= NOT \RegFile[13][13]~q\;
\ALT_INV_RegFile[30][29]~q\ <= NOT \RegFile[30][29]~q\;
\ALT_INV_RegFile[28][29]~q\ <= NOT \RegFile[28][29]~q\;
\ALT_INV_RegFile[31][29]~q\ <= NOT \RegFile[31][29]~q\;
\ALT_INV_RegFile[29][29]~q\ <= NOT \RegFile[29][29]~q\;
\ALT_INV_RegFile[22][29]~q\ <= NOT \RegFile[22][29]~q\;
\ALT_INV_RegFile[20][29]~q\ <= NOT \RegFile[20][29]~q\;
\ALT_INV_RegFile[23][29]~q\ <= NOT \RegFile[23][29]~q\;
\ALT_INV_RegFile[21][29]~q\ <= NOT \RegFile[21][29]~q\;
\ALT_INV_RegFile[14][29]~q\ <= NOT \RegFile[14][29]~q\;
\ALT_INV_RegFile[12][29]~q\ <= NOT \RegFile[12][29]~q\;
\ALT_INV_RegFile[15][29]~q\ <= NOT \RegFile[15][29]~q\;
\ALT_INV_RegFile[13][29]~q\ <= NOT \RegFile[13][29]~q\;
\ALT_INV_RegFile[30][4]~q\ <= NOT \RegFile[30][4]~q\;
\ALT_INV_RegFile[28][4]~q\ <= NOT \RegFile[28][4]~q\;
\ALT_INV_RegFile[31][4]~q\ <= NOT \RegFile[31][4]~q\;
\ALT_INV_RegFile[29][4]~q\ <= NOT \RegFile[29][4]~q\;
\ALT_INV_RegFile[22][4]~q\ <= NOT \RegFile[22][4]~q\;
\ALT_INV_RegFile[20][4]~q\ <= NOT \RegFile[20][4]~q\;
\ALT_INV_RegFile[23][4]~q\ <= NOT \RegFile[23][4]~q\;
\ALT_INV_RegFile[21][4]~q\ <= NOT \RegFile[21][4]~q\;
\ALT_INV_RegFile[14][4]~q\ <= NOT \RegFile[14][4]~q\;
\ALT_INV_RegFile[12][4]~q\ <= NOT \RegFile[12][4]~q\;
\ALT_INV_RegFile[15][4]~q\ <= NOT \RegFile[15][4]~q\;
\ALT_INV_RegFile[13][4]~q\ <= NOT \RegFile[13][4]~q\;
\ALT_INV_RegFile[30][12]~q\ <= NOT \RegFile[30][12]~q\;
\ALT_INV_RegFile[28][12]~q\ <= NOT \RegFile[28][12]~q\;
\ALT_INV_RegFile[31][12]~q\ <= NOT \RegFile[31][12]~q\;
\ALT_INV_RegFile[29][12]~q\ <= NOT \RegFile[29][12]~q\;
\ALT_INV_RegFile[22][12]~q\ <= NOT \RegFile[22][12]~q\;
\ALT_INV_RegFile[20][12]~q\ <= NOT \RegFile[20][12]~q\;
\ALT_INV_RegFile[23][12]~q\ <= NOT \RegFile[23][12]~q\;
\ALT_INV_RegFile[21][12]~q\ <= NOT \RegFile[21][12]~q\;
\ALT_INV_RegFile[14][12]~q\ <= NOT \RegFile[14][12]~q\;
\ALT_INV_RegFile[12][12]~q\ <= NOT \RegFile[12][12]~q\;
\ALT_INV_RegFile[15][12]~q\ <= NOT \RegFile[15][12]~q\;
\ALT_INV_RegFile[13][12]~q\ <= NOT \RegFile[13][12]~q\;
\ALT_INV_RegFile[30][28]~q\ <= NOT \RegFile[30][28]~q\;
\ALT_INV_RegFile[28][28]~q\ <= NOT \RegFile[28][28]~q\;
\ALT_INV_RegFile[31][28]~q\ <= NOT \RegFile[31][28]~q\;
\ALT_INV_RegFile[29][28]~q\ <= NOT \RegFile[29][28]~q\;
\ALT_INV_RegFile[22][28]~q\ <= NOT \RegFile[22][28]~q\;
\ALT_INV_RegFile[20][28]~q\ <= NOT \RegFile[20][28]~q\;
\ALT_INV_RegFile[23][28]~q\ <= NOT \RegFile[23][28]~q\;
\ALT_INV_RegFile[21][28]~q\ <= NOT \RegFile[21][28]~q\;
\ALT_INV_RegFile[14][28]~q\ <= NOT \RegFile[14][28]~q\;
\ALT_INV_RegFile[12][28]~q\ <= NOT \RegFile[12][28]~q\;
\ALT_INV_RegFile[15][28]~q\ <= NOT \RegFile[15][28]~q\;
\ALT_INV_RegFile[13][28]~q\ <= NOT \RegFile[13][28]~q\;
\ALT_INV_RegFile[30][3]~q\ <= NOT \RegFile[30][3]~q\;
\ALT_INV_RegFile[28][3]~q\ <= NOT \RegFile[28][3]~q\;
\ALT_INV_RegFile[31][3]~q\ <= NOT \RegFile[31][3]~q\;
\ALT_INV_RegFile[29][3]~q\ <= NOT \RegFile[29][3]~q\;
\ALT_INV_RegFile[22][3]~q\ <= NOT \RegFile[22][3]~q\;
\ALT_INV_RegFile[20][3]~q\ <= NOT \RegFile[20][3]~q\;
\ALT_INV_RegFile[23][3]~q\ <= NOT \RegFile[23][3]~q\;
\ALT_INV_RegFile[21][3]~q\ <= NOT \RegFile[21][3]~q\;
\ALT_INV_RegFile[14][3]~q\ <= NOT \RegFile[14][3]~q\;
\ALT_INV_RegFile[12][3]~q\ <= NOT \RegFile[12][3]~q\;
\ALT_INV_RegFile[15][3]~q\ <= NOT \RegFile[15][3]~q\;
\ALT_INV_RegFile[13][3]~q\ <= NOT \RegFile[13][3]~q\;
\ALT_INV_RegFile[30][11]~q\ <= NOT \RegFile[30][11]~q\;
\ALT_INV_RegFile[28][11]~q\ <= NOT \RegFile[28][11]~q\;
\ALT_INV_RegFile[31][11]~q\ <= NOT \RegFile[31][11]~q\;
\ALT_INV_RegFile[29][11]~q\ <= NOT \RegFile[29][11]~q\;
\ALT_INV_RegFile[22][11]~q\ <= NOT \RegFile[22][11]~q\;
\ALT_INV_RegFile[20][11]~q\ <= NOT \RegFile[20][11]~q\;
\ALT_INV_RegFile[23][11]~q\ <= NOT \RegFile[23][11]~q\;
\ALT_INV_RegFile[21][11]~q\ <= NOT \RegFile[21][11]~q\;
\ALT_INV_RegFile[14][11]~q\ <= NOT \RegFile[14][11]~q\;
\ALT_INV_RegFile[12][11]~q\ <= NOT \RegFile[12][11]~q\;
\ALT_INV_RegFile[15][11]~q\ <= NOT \RegFile[15][11]~q\;
\ALT_INV_RegFile[13][11]~q\ <= NOT \RegFile[13][11]~q\;
\ALT_INV_RegFile[30][27]~q\ <= NOT \RegFile[30][27]~q\;
\ALT_INV_RegFile[28][27]~q\ <= NOT \RegFile[28][27]~q\;
\ALT_INV_RegFile[31][27]~q\ <= NOT \RegFile[31][27]~q\;
\ALT_INV_RegFile[29][27]~q\ <= NOT \RegFile[29][27]~q\;
\ALT_INV_RegFile[22][27]~q\ <= NOT \RegFile[22][27]~q\;
\ALT_INV_RegFile[20][27]~q\ <= NOT \RegFile[20][27]~q\;
\ALT_INV_RegFile[23][27]~q\ <= NOT \RegFile[23][27]~q\;
\ALT_INV_RegFile[21][27]~q\ <= NOT \RegFile[21][27]~q\;
\ALT_INV_RegFile[14][27]~q\ <= NOT \RegFile[14][27]~q\;
\ALT_INV_RegFile[12][27]~q\ <= NOT \RegFile[12][27]~q\;
\ALT_INV_RegFile[15][27]~q\ <= NOT \RegFile[15][27]~q\;
\ALT_INV_RegFile[13][27]~q\ <= NOT \RegFile[13][27]~q\;
\ALT_INV_RegFile[30][2]~q\ <= NOT \RegFile[30][2]~q\;
\ALT_INV_RegFile[28][2]~q\ <= NOT \RegFile[28][2]~q\;
\ALT_INV_RegFile[31][2]~q\ <= NOT \RegFile[31][2]~q\;
\ALT_INV_RegFile[29][2]~q\ <= NOT \RegFile[29][2]~q\;
\ALT_INV_RegFile[22][2]~q\ <= NOT \RegFile[22][2]~q\;
\ALT_INV_RegFile[20][2]~q\ <= NOT \RegFile[20][2]~q\;
\ALT_INV_RegFile[23][2]~q\ <= NOT \RegFile[23][2]~q\;
\ALT_INV_RegFile[21][2]~q\ <= NOT \RegFile[21][2]~q\;
\ALT_INV_RegFile[14][2]~q\ <= NOT \RegFile[14][2]~q\;
\ALT_INV_RegFile[12][2]~q\ <= NOT \RegFile[12][2]~q\;
\ALT_INV_RegFile[15][2]~q\ <= NOT \RegFile[15][2]~q\;
\ALT_INV_RegFile[13][2]~q\ <= NOT \RegFile[13][2]~q\;
\ALT_INV_RegFile[30][10]~q\ <= NOT \RegFile[30][10]~q\;
\ALT_INV_RegFile[28][10]~q\ <= NOT \RegFile[28][10]~q\;
\ALT_INV_RegFile[31][10]~q\ <= NOT \RegFile[31][10]~q\;
\ALT_INV_RegFile[29][10]~q\ <= NOT \RegFile[29][10]~q\;
\ALT_INV_RegFile[22][10]~q\ <= NOT \RegFile[22][10]~q\;
\ALT_INV_RegFile[20][10]~q\ <= NOT \RegFile[20][10]~q\;
\ALT_INV_RegFile[23][10]~q\ <= NOT \RegFile[23][10]~q\;
\ALT_INV_RegFile[21][10]~q\ <= NOT \RegFile[21][10]~q\;
\ALT_INV_RegFile[14][10]~q\ <= NOT \RegFile[14][10]~q\;
\ALT_INV_RegFile[12][10]~q\ <= NOT \RegFile[12][10]~q\;
\ALT_INV_RegFile[15][10]~q\ <= NOT \RegFile[15][10]~q\;
\ALT_INV_RegFile[13][10]~q\ <= NOT \RegFile[13][10]~q\;
\ALT_INV_RegFile[30][26]~q\ <= NOT \RegFile[30][26]~q\;
\ALT_INV_RegFile[28][26]~q\ <= NOT \RegFile[28][26]~q\;
\ALT_INV_RegFile[31][26]~q\ <= NOT \RegFile[31][26]~q\;
\ALT_INV_RegFile[29][26]~q\ <= NOT \RegFile[29][26]~q\;
\ALT_INV_RegFile[22][26]~q\ <= NOT \RegFile[22][26]~q\;
\ALT_INV_RegFile[20][26]~q\ <= NOT \RegFile[20][26]~q\;
\ALT_INV_RegFile[23][26]~q\ <= NOT \RegFile[23][26]~q\;
\ALT_INV_RegFile[21][26]~q\ <= NOT \RegFile[21][26]~q\;
\ALT_INV_RegFile[14][26]~q\ <= NOT \RegFile[14][26]~q\;
\ALT_INV_RegFile[12][26]~q\ <= NOT \RegFile[12][26]~q\;
\ALT_INV_RegFile[15][26]~q\ <= NOT \RegFile[15][26]~q\;
\ALT_INV_RegFile[13][26]~q\ <= NOT \RegFile[13][26]~q\;
\ALT_INV_RegFile[30][1]~q\ <= NOT \RegFile[30][1]~q\;
\ALT_INV_RegFile[28][1]~q\ <= NOT \RegFile[28][1]~q\;
\ALT_INV_RegFile[31][1]~q\ <= NOT \RegFile[31][1]~q\;
\ALT_INV_RegFile[29][1]~q\ <= NOT \RegFile[29][1]~q\;
\ALT_INV_RegFile[22][1]~q\ <= NOT \RegFile[22][1]~q\;
\ALT_INV_RegFile[20][1]~q\ <= NOT \RegFile[20][1]~q\;
\ALT_INV_RegFile[23][1]~q\ <= NOT \RegFile[23][1]~q\;
\ALT_INV_RegFile[21][1]~q\ <= NOT \RegFile[21][1]~q\;
\ALT_INV_RegFile[14][1]~q\ <= NOT \RegFile[14][1]~q\;
\ALT_INV_RegFile[12][1]~q\ <= NOT \RegFile[12][1]~q\;
\ALT_INV_RegFile[15][1]~q\ <= NOT \RegFile[15][1]~q\;
\ALT_INV_RegFile[13][1]~q\ <= NOT \RegFile[13][1]~q\;
\ALT_INV_RegFile[30][9]~q\ <= NOT \RegFile[30][9]~q\;
\ALT_INV_RegFile[28][9]~q\ <= NOT \RegFile[28][9]~q\;
\ALT_INV_RegFile[31][9]~q\ <= NOT \RegFile[31][9]~q\;
\ALT_INV_RegFile[29][9]~q\ <= NOT \RegFile[29][9]~q\;
\ALT_INV_RegFile[22][9]~q\ <= NOT \RegFile[22][9]~q\;
\ALT_INV_RegFile[20][9]~q\ <= NOT \RegFile[20][9]~q\;
\ALT_INV_RegFile[23][9]~q\ <= NOT \RegFile[23][9]~q\;
\ALT_INV_RegFile[21][9]~q\ <= NOT \RegFile[21][9]~q\;
\ALT_INV_RegFile[14][9]~q\ <= NOT \RegFile[14][9]~q\;
\ALT_INV_RegFile[12][9]~q\ <= NOT \RegFile[12][9]~q\;
\ALT_INV_RegFile[15][9]~q\ <= NOT \RegFile[15][9]~q\;
\ALT_INV_RegFile[13][9]~q\ <= NOT \RegFile[13][9]~q\;
\ALT_INV_RegFile[30][25]~q\ <= NOT \RegFile[30][25]~q\;
\ALT_INV_RegFile[28][25]~q\ <= NOT \RegFile[28][25]~q\;
\ALT_INV_RegFile[31][25]~q\ <= NOT \RegFile[31][25]~q\;
\ALT_INV_RegFile[29][25]~q\ <= NOT \RegFile[29][25]~q\;
\ALT_INV_RegFile[22][25]~q\ <= NOT \RegFile[22][25]~q\;
\ALT_INV_RegFile[20][25]~q\ <= NOT \RegFile[20][25]~q\;
\ALT_INV_RegFile[23][25]~q\ <= NOT \RegFile[23][25]~q\;
\ALT_INV_RegFile[21][25]~q\ <= NOT \RegFile[21][25]~q\;
\ALT_INV_RegFile[14][25]~q\ <= NOT \RegFile[14][25]~q\;
\ALT_INV_RegFile[12][25]~q\ <= NOT \RegFile[12][25]~q\;
\ALT_INV_RegFile[15][25]~q\ <= NOT \RegFile[15][25]~q\;
\ALT_INV_RegFile[13][25]~q\ <= NOT \RegFile[13][25]~q\;
\ALT_INV_RegFile[30][0]~q\ <= NOT \RegFile[30][0]~q\;
\ALT_INV_RegFile[28][0]~q\ <= NOT \RegFile[28][0]~q\;
\ALT_INV_RegFile[31][0]~q\ <= NOT \RegFile[31][0]~q\;
\ALT_INV_RegFile[29][0]~q\ <= NOT \RegFile[29][0]~q\;
\ALT_INV_RegFile[22][0]~q\ <= NOT \RegFile[22][0]~q\;
\ALT_INV_RegFile[20][0]~q\ <= NOT \RegFile[20][0]~q\;
\ALT_INV_RegFile[23][0]~q\ <= NOT \RegFile[23][0]~q\;
\ALT_INV_RegFile[21][0]~q\ <= NOT \RegFile[21][0]~q\;
\ALT_INV_RegFile[14][0]~q\ <= NOT \RegFile[14][0]~q\;
\ALT_INV_RegFile[12][0]~q\ <= NOT \RegFile[12][0]~q\;
\ALT_INV_RegFile[15][0]~q\ <= NOT \RegFile[15][0]~q\;
\ALT_INV_RegFile[13][0]~q\ <= NOT \RegFile[13][0]~q\;
\ALT_INV_RegFile[30][8]~q\ <= NOT \RegFile[30][8]~q\;
\ALT_INV_RegFile[28][8]~q\ <= NOT \RegFile[28][8]~q\;
\ALT_INV_RegFile[31][8]~q\ <= NOT \RegFile[31][8]~q\;
\ALT_INV_RegFile[29][8]~q\ <= NOT \RegFile[29][8]~q\;
\ALT_INV_RegFile[22][8]~q\ <= NOT \RegFile[22][8]~q\;
\ALT_INV_RegFile[20][8]~q\ <= NOT \RegFile[20][8]~q\;
\ALT_INV_RegFile[23][8]~q\ <= NOT \RegFile[23][8]~q\;
\ALT_INV_RegFile[21][8]~q\ <= NOT \RegFile[21][8]~q\;
\ALT_INV_RegFile[14][8]~q\ <= NOT \RegFile[14][8]~q\;
\ALT_INV_RegFile[12][8]~q\ <= NOT \RegFile[12][8]~q\;
\ALT_INV_RegFile[15][8]~q\ <= NOT \RegFile[15][8]~q\;
\ALT_INV_RegFile[13][8]~q\ <= NOT \RegFile[13][8]~q\;
\ALT_INV_RegFile[30][24]~q\ <= NOT \RegFile[30][24]~q\;
\ALT_INV_RegFile[28][24]~q\ <= NOT \RegFile[28][24]~q\;
\ALT_INV_RegFile[31][24]~q\ <= NOT \RegFile[31][24]~q\;
\ALT_INV_RegFile[29][24]~q\ <= NOT \RegFile[29][24]~q\;
\ALT_INV_RegFile[22][24]~q\ <= NOT \RegFile[22][24]~q\;
\ALT_INV_RegFile[20][24]~q\ <= NOT \RegFile[20][24]~q\;
\ALT_INV_RegFile[23][24]~q\ <= NOT \RegFile[23][24]~q\;
\ALT_INV_RegFile[21][24]~q\ <= NOT \RegFile[21][24]~q\;
\ALT_INV_RegFile[14][24]~q\ <= NOT \RegFile[14][24]~q\;
\ALT_INV_RegFile[12][24]~q\ <= NOT \RegFile[12][24]~q\;
\ALT_INV_RegFile[15][24]~q\ <= NOT \RegFile[15][24]~q\;
\ALT_INV_RegFile[13][24]~q\ <= NOT \RegFile[13][24]~q\;
\ALT_INV_R.regWriteEn~q\ <= NOT \R.regWriteEn~q\;
\ALT_INV_Selector23~6_combout\ <= NOT \Selector23~6_combout\;
\ALT_INV_Selector25~6_combout\ <= NOT \Selector25~6_combout\;
\ALT_INV_Mux21~2_combout\ <= NOT \Mux21~2_combout\;
\ALT_INV_Mux21~1_combout\ <= NOT \Mux21~1_combout\;
\ALT_INV_Mux22~1_combout\ <= NOT \Mux22~1_combout\;
\ALT_INV_Mux22~0_combout\ <= NOT \Mux22~0_combout\;
\ALT_INV_Mux24~1_combout\ <= NOT \Mux24~1_combout\;
\ALT_INV_Mux24~0_combout\ <= NOT \Mux24~0_combout\;
\ALT_INV_Mux18~1_combout\ <= NOT \Mux18~1_combout\;
\ALT_INV_Mux17~1_combout\ <= NOT \Mux17~1_combout\;
\ALT_INV_Mux17~0_combout\ <= NOT \Mux17~0_combout\;
\ALT_INV_Comb~1_combout\ <= NOT \Comb~1_combout\;
\ALT_INV_Mux0~0_combout\ <= NOT \Mux0~0_combout\;
\ALT_INV_Mux23~1_combout\ <= NOT \Mux23~1_combout\;
\ALT_INV_Mux23~0_combout\ <= NOT \Mux23~0_combout\;
\ALT_INV_Mux26~2_combout\ <= NOT \Mux26~2_combout\;
\ALT_INV_Mux26~1_combout\ <= NOT \Mux26~1_combout\;
\ALT_INV_Mux25~1_combout\ <= NOT \Mux25~1_combout\;
\ALT_INV_Mux25~0_combout\ <= NOT \Mux25~0_combout\;
\ALT_INV_Mux21~0_combout\ <= NOT \Mux21~0_combout\;
\ALT_INV_Mux125~0_combout\ <= NOT \Mux125~0_combout\;
\ALT_INV_Mux225~0_combout\ <= NOT \Mux225~0_combout\;
\ALT_INV_Mux61~13_combout\ <= NOT \Mux61~13_combout\;
\ALT_INV_Mux61~0_combout\ <= NOT \Mux61~0_combout\;
\ALT_INV_Mux124~1_combout\ <= NOT \Mux124~1_combout\;
\ALT_INV_Mux224~0_combout\ <= NOT \Mux224~0_combout\;
\ALT_INV_Mux60~13_combout\ <= NOT \Mux60~13_combout\;
\ALT_INV_Mux60~0_combout\ <= NOT \Mux60~0_combout\;
\ALT_INV_NxR.aluData2[31]~29_combout\ <= NOT \NxR.aluData2[31]~29_combout\;
\ALT_INV_Mux123~3_combout\ <= NOT \Mux123~3_combout\;
\ALT_INV_Mux223~0_combout\ <= NOT \Mux223~0_combout\;
\ALT_INV_Mux59~13_combout\ <= NOT \Mux59~13_combout\;
\ALT_INV_Mux59~0_combout\ <= NOT \Mux59~0_combout\;
\ALT_INV_Mux132~0_combout\ <= NOT \Mux132~0_combout\;
\ALT_INV_Mux232~0_combout\ <= NOT \Mux232~0_combout\;
\ALT_INV_Mux68~13_combout\ <= NOT \Mux68~13_combout\;
\ALT_INV_Mux68~0_combout\ <= NOT \Mux68~0_combout\;
\ALT_INV_Mux131~0_combout\ <= NOT \Mux131~0_combout\;
\ALT_INV_Mux231~0_combout\ <= NOT \Mux231~0_combout\;
\ALT_INV_Mux67~13_combout\ <= NOT \Mux67~13_combout\;
\ALT_INV_Mux67~0_combout\ <= NOT \Mux67~0_combout\;
\ALT_INV_Mux130~0_combout\ <= NOT \Mux130~0_combout\;
\ALT_INV_Mux230~0_combout\ <= NOT \Mux230~0_combout\;
\ALT_INV_Mux66~13_combout\ <= NOT \Mux66~13_combout\;
\ALT_INV_Mux66~0_combout\ <= NOT \Mux66~0_combout\;
\ALT_INV_NxR.aluData2[26]~25_combout\ <= NOT \NxR.aluData2[26]~25_combout\;
\ALT_INV_Mux128~0_combout\ <= NOT \Mux128~0_combout\;
\ALT_INV_Mux228~0_combout\ <= NOT \Mux228~0_combout\;
\ALT_INV_Mux64~13_combout\ <= NOT \Mux64~13_combout\;
\ALT_INV_Mux64~0_combout\ <= NOT \Mux64~0_combout\;
\ALT_INV_NxR.aluData2[27]~24_combout\ <= NOT \NxR.aluData2[27]~24_combout\;
\ALT_INV_Mux127~0_combout\ <= NOT \Mux127~0_combout\;
\ALT_INV_Mux227~0_combout\ <= NOT \Mux227~0_combout\;
\ALT_INV_Mux63~13_combout\ <= NOT \Mux63~13_combout\;
\ALT_INV_Mux63~0_combout\ <= NOT \Mux63~0_combout\;
\ALT_INV_NxR.aluData2[28]~23_combout\ <= NOT \NxR.aluData2[28]~23_combout\;
\ALT_INV_Mux126~0_combout\ <= NOT \Mux126~0_combout\;
\ALT_INV_Mux226~0_combout\ <= NOT \Mux226~0_combout\;
\ALT_INV_Mux62~13_combout\ <= NOT \Mux62~13_combout\;
\ALT_INV_Mux62~0_combout\ <= NOT \Mux62~0_combout\;
\ALT_INV_Mux129~0_combout\ <= NOT \Mux129~0_combout\;
\ALT_INV_Mux229~0_combout\ <= NOT \Mux229~0_combout\;
\ALT_INV_Mux65~13_combout\ <= NOT \Mux65~13_combout\;
\ALT_INV_Mux65~0_combout\ <= NOT \Mux65~0_combout\;
\ALT_INV_Mux250~0_combout\ <= NOT \Mux250~0_combout\;
\ALT_INV_Mux86~13_combout\ <= NOT \Mux86~13_combout\;
\ALT_INV_Mux86~0_combout\ <= NOT \Mux86~0_combout\;
\ALT_INV_NxR.aluData2[5]~21_combout\ <= NOT \NxR.aluData2[5]~21_combout\;
\ALT_INV_Mux149~1_combout\ <= NOT \Mux149~1_combout\;
\ALT_INV_Mux249~0_combout\ <= NOT \Mux249~0_combout\;
\ALT_INV_Mux85~13_combout\ <= NOT \Mux85~13_combout\;
\ALT_INV_Mux85~0_combout\ <= NOT \Mux85~0_combout\;
\ALT_INV_NxR.aluData2[4]~20_combout\ <= NOT \NxR.aluData2[4]~20_combout\;
\ALT_INV_Mux150~0_combout\ <= NOT \Mux150~0_combout\;
\ALT_INV_R.curInst\(11) <= NOT \R.curInst\(11);
\ALT_INV_Mux252~0_combout\ <= NOT \Mux252~0_combout\;
\ALT_INV_Mux88~13_combout\ <= NOT \Mux88~13_combout\;
\ALT_INV_Mux88~0_combout\ <= NOT \Mux88~0_combout\;
\ALT_INV_Mux251~0_combout\ <= NOT \Mux251~0_combout\;
\ALT_INV_Mux87~13_combout\ <= NOT \Mux87~13_combout\;
\ALT_INV_Mux87~0_combout\ <= NOT \Mux87~0_combout\;
\ALT_INV_NxR.aluData2[2]~19_combout\ <= NOT \NxR.aluData2[2]~19_combout\;
\ALT_INV_Mux152~0_combout\ <= NOT \Mux152~0_combout\;
\ALT_INV_R.curInst\(9) <= NOT \R.curInst\(9);
\ALT_INV_NxR.aluData2[3]~18_combout\ <= NOT \NxR.aluData2[3]~18_combout\;
\ALT_INV_Mux151~0_combout\ <= NOT \Mux151~0_combout\;
\ALT_INV_R.curInst\(10) <= NOT \R.curInst\(10);
\ALT_INV_Mux253~0_combout\ <= NOT \Mux253~0_combout\;
\ALT_INV_Mux89~13_combout\ <= NOT \Mux89~13_combout\;
\ALT_INV_Mux89~0_combout\ <= NOT \Mux89~0_combout\;
\ALT_INV_NxR.aluData2[1]~17_combout\ <= NOT \NxR.aluData2[1]~17_combout\;
\ALT_INV_Mux153~0_combout\ <= NOT \Mux153~0_combout\;
\ALT_INV_R.curInst\(8) <= NOT \R.curInst\(8);
\ALT_INV_NxR.aluData2[0]~16_combout\ <= NOT \NxR.aluData2[0]~16_combout\;
\ALT_INV_Mux154~1_combout\ <= NOT \Mux154~1_combout\;
\ALT_INV_Mux254~0_combout\ <= NOT \Mux254~0_combout\;
\ALT_INV_Mux90~13_combout\ <= NOT \Mux90~13_combout\;
\ALT_INV_Mux90~0_combout\ <= NOT \Mux90~0_combout\;
\ALT_INV_NxR.aluData2[6]~15_combout\ <= NOT \NxR.aluData2[6]~15_combout\;
\ALT_INV_Mux148~0_combout\ <= NOT \Mux148~0_combout\;
\ALT_INV_Mux248~0_combout\ <= NOT \Mux248~0_combout\;
\ALT_INV_Mux84~13_combout\ <= NOT \Mux84~13_combout\;
\ALT_INV_Mux84~0_combout\ <= NOT \Mux84~0_combout\;
\ALT_INV_NxR.aluData2[7]~14_combout\ <= NOT \NxR.aluData2[7]~14_combout\;
\ALT_INV_Mux147~0_combout\ <= NOT \Mux147~0_combout\;
\ALT_INV_Mux247~0_combout\ <= NOT \Mux247~0_combout\;
\ALT_INV_Mux83~13_combout\ <= NOT \Mux83~13_combout\;
\ALT_INV_Mux83~0_combout\ <= NOT \Mux83~0_combout\;
\ALT_INV_NxR.aluData2[8]~13_combout\ <= NOT \NxR.aluData2[8]~13_combout\;
\ALT_INV_Mux146~0_combout\ <= NOT \Mux146~0_combout\;
\ALT_INV_Mux246~0_combout\ <= NOT \Mux246~0_combout\;
\ALT_INV_Mux82~13_combout\ <= NOT \Mux82~13_combout\;
\ALT_INV_Mux82~0_combout\ <= NOT \Mux82~0_combout\;
\ALT_INV_NxR.aluData2[9]~12_combout\ <= NOT \NxR.aluData2[9]~12_combout\;
\ALT_INV_Mux145~0_combout\ <= NOT \Mux145~0_combout\;
\ALT_INV_Mux245~0_combout\ <= NOT \Mux245~0_combout\;
\ALT_INV_Mux81~13_combout\ <= NOT \Mux81~13_combout\;
\ALT_INV_Mux81~0_combout\ <= NOT \Mux81~0_combout\;
\ALT_INV_NxR.aluData2[12]~11_combout\ <= NOT \NxR.aluData2[12]~11_combout\;
\ALT_INV_Mux142~0_combout\ <= NOT \Mux142~0_combout\;
\ALT_INV_Mux242~0_combout\ <= NOT \Mux242~0_combout\;
\ALT_INV_Mux78~13_combout\ <= NOT \Mux78~13_combout\;
\ALT_INV_Mux78~0_combout\ <= NOT \Mux78~0_combout\;
\ALT_INV_NxR.aluData2[13]~10_combout\ <= NOT \NxR.aluData2[13]~10_combout\;
\ALT_INV_Mux141~0_combout\ <= NOT \Mux141~0_combout\;
\ALT_INV_Mux241~0_combout\ <= NOT \Mux241~0_combout\;
\ALT_INV_Mux77~13_combout\ <= NOT \Mux77~13_combout\;
\ALT_INV_Mux77~0_combout\ <= NOT \Mux77~0_combout\;
\ALT_INV_NxR.aluData2[10]~9_combout\ <= NOT \NxR.aluData2[10]~9_combout\;
\ALT_INV_Mux144~0_combout\ <= NOT \Mux144~0_combout\;
\ALT_INV_Mux244~0_combout\ <= NOT \Mux244~0_combout\;
\ALT_INV_Mux80~13_combout\ <= NOT \Mux80~13_combout\;
\ALT_INV_Mux80~0_combout\ <= NOT \Mux80~0_combout\;
\ALT_INV_NxR.aluData2[11]~8_combout\ <= NOT \NxR.aluData2[11]~8_combout\;
\ALT_INV_Mux143~1_combout\ <= NOT \Mux143~1_combout\;
\ALT_INV_Mux143~0_combout\ <= NOT \Mux143~0_combout\;
\ALT_INV_R.curInst\(7) <= NOT \R.curInst\(7);
\ALT_INV_Mux243~0_combout\ <= NOT \Mux243~0_combout\;
\ALT_INV_Mux79~13_combout\ <= NOT \Mux79~13_combout\;
\ALT_INV_Mux79~0_combout\ <= NOT \Mux79~0_combout\;
\ALT_INV_NxR.aluData2[14]~7_combout\ <= NOT \NxR.aluData2[14]~7_combout\;
\ALT_INV_Mux140~0_combout\ <= NOT \Mux140~0_combout\;

-- Location: IOOBUF_X40_Y81_N2
\avm_i_address[0]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC[0]~DUPLICATE_q\,
	devoe => ww_devoe,
	o => ww_avm_i_address(0));

-- Location: IOOBUF_X22_Y0_N19
\avm_i_address[1]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(1),
	devoe => ww_devoe,
	o => ww_avm_i_address(1));

-- Location: IOOBUF_X89_Y15_N22
\avm_i_address[2]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(2),
	devoe => ww_devoe,
	o => ww_avm_i_address(2));

-- Location: IOOBUF_X89_Y16_N5
\avm_i_address[3]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(3),
	devoe => ww_devoe,
	o => ww_avm_i_address(3));

-- Location: IOOBUF_X89_Y15_N39
\avm_i_address[4]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(4),
	devoe => ww_devoe,
	o => ww_avm_i_address(4));

-- Location: IOOBUF_X89_Y11_N79
\avm_i_address[5]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(5),
	devoe => ww_devoe,
	o => ww_avm_i_address(5));

-- Location: IOOBUF_X89_Y15_N5
\avm_i_address[6]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(6),
	devoe => ww_devoe,
	o => ww_avm_i_address(6));

-- Location: IOOBUF_X89_Y13_N56
\avm_i_address[7]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(7),
	devoe => ww_devoe,
	o => ww_avm_i_address(7));

-- Location: IOOBUF_X89_Y13_N5
\avm_i_address[8]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(8),
	devoe => ww_devoe,
	o => ww_avm_i_address(8));

-- Location: IOOBUF_X86_Y0_N19
\avm_i_address[9]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(9),
	devoe => ww_devoe,
	o => ww_avm_i_address(9));

-- Location: IOOBUF_X89_Y8_N39
\avm_i_address[10]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(10),
	devoe => ww_devoe,
	o => ww_avm_i_address(10));

-- Location: IOOBUF_X89_Y6_N22
\avm_i_address[11]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(11),
	devoe => ww_devoe,
	o => ww_avm_i_address(11));

-- Location: IOOBUF_X89_Y8_N5
\avm_i_address[12]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(12),
	devoe => ww_devoe,
	o => ww_avm_i_address(12));

-- Location: IOOBUF_X89_Y11_N96
\avm_i_address[13]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(13),
	devoe => ww_devoe,
	o => ww_avm_i_address(13));

-- Location: IOOBUF_X89_Y6_N39
\avm_i_address[14]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(14),
	devoe => ww_devoe,
	o => ww_avm_i_address(14));

-- Location: IOOBUF_X89_Y6_N56
\avm_i_address[15]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(15),
	devoe => ww_devoe,
	o => ww_avm_i_address(15));

-- Location: IOOBUF_X89_Y4_N79
\avm_i_address[16]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(16),
	devoe => ww_devoe,
	o => ww_avm_i_address(16));

-- Location: IOOBUF_X62_Y0_N36
\avm_i_address[17]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(17),
	devoe => ww_devoe,
	o => ww_avm_i_address(17));

-- Location: IOOBUF_X70_Y0_N19
\avm_i_address[18]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(18),
	devoe => ww_devoe,
	o => ww_avm_i_address(18));

-- Location: IOOBUF_X89_Y6_N5
\avm_i_address[19]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(19),
	devoe => ww_devoe,
	o => ww_avm_i_address(19));

-- Location: IOOBUF_X89_Y8_N22
\avm_i_address[20]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(20),
	devoe => ww_devoe,
	o => ww_avm_i_address(20));

-- Location: IOOBUF_X62_Y0_N2
\avm_i_address[21]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC[21]~DUPLICATE_q\,
	devoe => ww_devoe,
	o => ww_avm_i_address(21));

-- Location: IOOBUF_X82_Y0_N59
\avm_i_address[22]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(22),
	devoe => ww_devoe,
	o => ww_avm_i_address(22));

-- Location: IOOBUF_X89_Y4_N96
\avm_i_address[23]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(23),
	devoe => ww_devoe,
	o => ww_avm_i_address(23));

-- Location: IOOBUF_X89_Y4_N62
\avm_i_address[24]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(24),
	devoe => ww_devoe,
	o => ww_avm_i_address(24));

-- Location: IOOBUF_X82_Y0_N42
\avm_i_address[25]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(25),
	devoe => ww_devoe,
	o => ww_avm_i_address(25));

-- Location: IOOBUF_X70_Y0_N2
\avm_i_address[26]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(26),
	devoe => ww_devoe,
	o => ww_avm_i_address(26));

-- Location: IOOBUF_X82_Y0_N76
\avm_i_address[27]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(27),
	devoe => ww_devoe,
	o => ww_avm_i_address(27));

-- Location: IOOBUF_X72_Y0_N53
\avm_i_address[28]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC\(28),
	devoe => ww_devoe,
	o => ww_avm_i_address(28));

-- Location: IOOBUF_X88_Y0_N54
\avm_i_address[29]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC[29]~DUPLICATE_q\,
	devoe => ww_devoe,
	o => ww_avm_i_address(29));

-- Location: IOOBUF_X32_Y0_N2
\avm_i_address[30]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC[30]~DUPLICATE_q\,
	devoe => ww_devoe,
	o => ww_avm_i_address(30));

-- Location: IOOBUF_X26_Y0_N59
\avm_i_address[31]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.curPC[31]~DUPLICATE_q\,
	devoe => ww_devoe,
	o => ww_avm_i_address(31));

-- Location: IOOBUF_X58_Y0_N42
\avm_i_read~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Comb~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_i_read);

-- Location: IOOBUF_X89_Y16_N39
\avm_d_address[0]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(0));

-- Location: IOOBUF_X89_Y13_N39
\avm_d_address[1]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~1_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(1));

-- Location: IOOBUF_X89_Y11_N45
\avm_d_address[2]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~2_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(2));

-- Location: IOOBUF_X89_Y9_N5
\avm_d_address[3]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~3_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(3));

-- Location: IOOBUF_X38_Y81_N36
\avm_d_address[4]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~4_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(4));

-- Location: IOOBUF_X89_Y8_N56
\avm_d_address[5]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~5_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(5));

-- Location: IOOBUF_X89_Y9_N22
\avm_d_address[6]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~6_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(6));

-- Location: IOOBUF_X89_Y9_N39
\avm_d_address[7]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~7_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(7));

-- Location: IOOBUF_X38_Y81_N2
\avm_d_address[8]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~8_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(8));

-- Location: IOOBUF_X32_Y0_N36
\avm_d_address[9]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~9_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(9));

-- Location: IOOBUF_X89_Y20_N96
\avm_d_address[10]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~10_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(10));

-- Location: IOOBUF_X89_Y16_N22
\avm_d_address[11]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~60_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(11));

-- Location: IOOBUF_X38_Y81_N53
\avm_d_address[12]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~11_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(12));

-- Location: IOOBUF_X89_Y15_N56
\avm_d_address[13]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~56_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(13));

-- Location: IOOBUF_X24_Y0_N53
\avm_d_address[14]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~12_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(14));

-- Location: IOOBUF_X89_Y21_N5
\avm_d_address[15]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~52_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(15));

-- Location: IOOBUF_X38_Y0_N36
\avm_d_address[16]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~13_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(16));

-- Location: IOOBUF_X30_Y0_N19
\avm_d_address[17]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~14_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(17));

-- Location: IOOBUF_X30_Y0_N2
\avm_d_address[18]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~15_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(18));

-- Location: IOOBUF_X86_Y0_N53
\avm_d_address[19]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~16_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(19));

-- Location: IOOBUF_X89_Y20_N62
\avm_d_address[20]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~17_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(20));

-- Location: IOOBUF_X58_Y0_N59
\avm_d_address[21]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~18_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(21));

-- Location: IOOBUF_X60_Y0_N36
\avm_d_address[22]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~19_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(22));

-- Location: IOOBUF_X86_Y0_N2
\avm_d_address[23]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~20_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(23));

-- Location: IOOBUF_X86_Y0_N36
\avm_d_address[24]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~21_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(24));

-- Location: IOOBUF_X89_Y9_N56
\avm_d_address[25]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~22_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(25));

-- Location: IOOBUF_X24_Y0_N36
\avm_d_address[26]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~23_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(26));

-- Location: IOOBUF_X89_Y20_N79
\avm_d_address[27]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~24_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(27));

-- Location: IOOBUF_X26_Y0_N42
\avm_d_address[28]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~48_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(28));

-- Location: IOOBUF_X88_Y0_N3
\avm_d_address[29]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~44_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(29));

-- Location: IOOBUF_X34_Y81_N42
\avm_d_address[30]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~40_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(30));

-- Location: IOOBUF_X40_Y81_N36
\avm_d_address[31]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \vAluRes~36_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_address(31));

-- Location: IOOBUF_X88_Y0_N37
\avm_d_byteenable[0]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux222~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_byteenable(0));

-- Location: IOOBUF_X50_Y0_N93
\avm_d_byteenable[1]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux221~1_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_byteenable(1));

-- Location: IOOBUF_X28_Y0_N53
\avm_d_byteenable[2]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux221~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_byteenable(2));

-- Location: IOOBUF_X28_Y0_N2
\avm_d_byteenable[3]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux221~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_byteenable(3));

-- Location: IOOBUF_X32_Y0_N53
\avm_d_write~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.memWrite~q\,
	devoe => ww_devoe,
	o => ww_avm_d_write);

-- Location: IOOBUF_X56_Y0_N36
\avm_d_writedata[0]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux194~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(0));

-- Location: IOOBUF_X54_Y0_N2
\avm_d_writedata[1]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux193~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(1));

-- Location: IOOBUF_X54_Y0_N19
\avm_d_writedata[2]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux192~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(2));

-- Location: IOOBUF_X30_Y0_N36
\avm_d_writedata[3]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux191~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(3));

-- Location: IOOBUF_X28_Y0_N36
\avm_d_writedata[4]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux190~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(4));

-- Location: IOOBUF_X54_Y0_N36
\avm_d_writedata[5]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux189~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(5));

-- Location: IOOBUF_X36_Y0_N36
\avm_d_writedata[6]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux188~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(6));

-- Location: IOOBUF_X30_Y0_N53
\avm_d_writedata[7]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux187~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(7));

-- Location: IOOBUF_X60_Y0_N19
\avm_d_writedata[8]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux202~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(8));

-- Location: IOOBUF_X52_Y0_N19
\avm_d_writedata[9]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux201~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(9));

-- Location: IOOBUF_X56_Y0_N2
\avm_d_writedata[10]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux200~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(10));

-- Location: IOOBUF_X38_Y81_N19
\avm_d_writedata[11]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux199~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(11));

-- Location: IOOBUF_X52_Y0_N2
\avm_d_writedata[12]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux198~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(12));

-- Location: IOOBUF_X50_Y0_N59
\avm_d_writedata[13]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux197~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(13));

-- Location: IOOBUF_X52_Y0_N36
\avm_d_writedata[14]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux196~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(14));

-- Location: IOOBUF_X56_Y0_N19
\avm_d_writedata[15]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux195~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(15));

-- Location: IOOBUF_X16_Y0_N36
\avm_d_writedata[16]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux210~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(16));

-- Location: IOOBUF_X38_Y0_N19
\avm_d_writedata[17]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux209~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(17));

-- Location: IOOBUF_X38_Y0_N2
\avm_d_writedata[18]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux208~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(18));

-- Location: IOOBUF_X28_Y0_N19
\avm_d_writedata[19]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux207~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(19));

-- Location: IOOBUF_X40_Y0_N53
\avm_d_writedata[20]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux206~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(20));

-- Location: IOOBUF_X50_Y0_N42
\avm_d_writedata[21]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux205~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(21));

-- Location: IOOBUF_X40_Y0_N2
\avm_d_writedata[22]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux204~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(22));

-- Location: IOOBUF_X52_Y0_N53
\avm_d_writedata[23]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux203~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(23));

-- Location: IOOBUF_X50_Y0_N76
\avm_d_writedata[24]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux218~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(24));

-- Location: IOOBUF_X89_Y4_N45
\avm_d_writedata[25]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux217~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(25));

-- Location: IOOBUF_X89_Y16_N56
\avm_d_writedata[26]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux216~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(26));

-- Location: IOOBUF_X40_Y0_N36
\avm_d_writedata[27]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux215~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(27));

-- Location: IOOBUF_X38_Y0_N53
\avm_d_writedata[28]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux214~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(28));

-- Location: IOOBUF_X40_Y81_N53
\avm_d_writedata[29]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux213~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(29));

-- Location: IOOBUF_X40_Y0_N19
\avm_d_writedata[30]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux212~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(30));

-- Location: IOOBUF_X40_Y81_N19
\avm_d_writedata[31]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Mux211~0_combout\,
	devoe => ww_devoe,
	o => ww_avm_d_writedata(31));

-- Location: IOOBUF_X34_Y0_N42
\avm_d_read~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \R.memRead~q\,
	devoe => ww_devoe,
	o => ww_avm_d_read);

-- Location: IOIBUF_X89_Y25_N21
\csi_clk~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_csi_clk,
	o => \csi_clk~input_o\);

-- Location: CLKCTRL_G10
\csi_clk~inputCLKENA0\ : cyclonev_clkena
-- pragma translate_off
GENERIC MAP (
	clock_type => "global clock",
	disable_mode => "low",
	ena_register_mode => "always enabled",
	ena_register_power_up => "high",
	test_syn => "high")
-- pragma translate_on
PORT MAP (
	inclk => \csi_clk~input_o\,
	outclk => \csi_clk~inputCLKENA0_outclk\);

-- Location: IOIBUF_X72_Y0_N18
\avm_i_readdata[31]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(31),
	o => \avm_i_readdata[31]~input_o\);

-- Location: IOIBUF_X89_Y23_N4
\rsi_reset_n~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_rsi_reset_n,
	o => \rsi_reset_n~input_o\);

-- Location: CLKCTRL_G8
\rsi_reset_n~inputCLKENA0\ : cyclonev_clkena
-- pragma translate_off
GENERIC MAP (
	clock_type => "global clock",
	disable_mode => "low",
	ena_register_mode => "always enabled",
	ena_register_power_up => "high",
	test_syn => "high")
-- pragma translate_on
PORT MAP (
	inclk => \rsi_reset_n~input_o\,
	outclk => \rsi_reset_n~inputCLKENA0_outclk\);

-- Location: DDIOINCELL_X72_Y0_N31
\R.curInst[7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[31]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(7));

-- Location: IOIBUF_X76_Y0_N18
\avm_i_readdata[26]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(26),
	o => \avm_i_readdata[26]~input_o\);

-- Location: DDIOINCELL_X76_Y0_N31
\R.curInst[2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[26]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(2));

-- Location: IOIBUF_X76_Y0_N35
\avm_i_readdata[28]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(28),
	o => \avm_i_readdata[28]~input_o\);

-- Location: DDIOINCELL_X76_Y0_N48
\R.curInst[4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[28]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(4));

-- Location: IOIBUF_X76_Y0_N1
\avm_i_readdata[30]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(30),
	o => \avm_i_readdata[30]~input_o\);

-- Location: DDIOINCELL_X76_Y0_N14
\R.curInst[6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[30]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(6));

-- Location: IOIBUF_X76_Y0_N52
\avm_i_readdata[29]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(29),
	o => \avm_i_readdata[29]~input_o\);

-- Location: DDIOINCELL_X76_Y0_N65
\R.curInst[5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[29]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(5));

-- Location: IOIBUF_X66_Y0_N75
\avm_i_readdata[12]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(12),
	o => \avm_i_readdata[12]~input_o\);

-- Location: DDIOINCELL_X66_Y0_N88
\R.curInst[20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[12]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(20));

-- Location: LABCELL_X77_Y2_N54
\Mux154~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux154~1_combout\ = ( \R.curInst\(5) & ( \R.curInst\(20) & ( (!\R.curInst\(4) & ((!\R.curInst\(2) & (\R.curInst\(7) & !\R.curInst\(6))) # (\R.curInst\(2) & ((\R.curInst\(6)))))) ) ) ) # ( !\R.curInst\(5) & ( \R.curInst\(20) & ( (!\R.curInst\(2) & 
-- !\R.curInst\(6)) ) ) ) # ( \R.curInst\(5) & ( !\R.curInst\(20) & ( (\R.curInst\(7) & (!\R.curInst\(2) & (!\R.curInst\(4) & !\R.curInst\(6)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010000000000000011001100000000000100000000110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(7),
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_R.curInst\(4),
	datad => \ALT_INV_R.curInst\(6),
	datae => \ALT_INV_R.curInst\(5),
	dataf => \ALT_INV_R.curInst\(20),
	combout => \Mux154~1_combout\);

-- Location: IOIBUF_X78_Y0_N52
\avm_i_readdata[27]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(27),
	o => \avm_i_readdata[27]~input_o\);

-- Location: DDIOINCELL_X78_Y0_N65
\R.curInst[3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[27]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(3));

-- Location: IOIBUF_X78_Y0_N35
\avm_i_readdata[24]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(24),
	o => \avm_i_readdata[24]~input_o\);

-- Location: DDIOINCELL_X78_Y0_N48
\R.curInst[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[24]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(0));

-- Location: IOIBUF_X78_Y0_N1
\avm_i_readdata[25]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(25),
	o => \avm_i_readdata[25]~input_o\);

-- Location: DDIOINCELL_X78_Y0_N14
\R.curInst[1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[25]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(1));

-- Location: LABCELL_X74_Y4_N12
\Equal4~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Equal4~1_combout\ = ( \R.curInst\(1) & ( \R.curInst\(0) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000111111110000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \ALT_INV_R.curInst\(0),
	dataf => \ALT_INV_R.curInst\(1),
	combout => \Equal4~1_combout\);

-- Location: LABCELL_X77_Y1_N57
\Mux34~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux34~0_combout\ = ( \R.curInst\(6) & ( \R.curInst\(5) & ( (!\R.curInst\(2) & (!\R.curInst\(3))) # (\R.curInst\(2) & ((!\R.curInst\(4)))) ) ) ) # ( !\R.curInst\(6) & ( \R.curInst\(5) & ( (!\R.curInst\(3) & ((!\R.curInst\(2)) # (\R.curInst\(4)))) ) ) ) # 
-- ( !\R.curInst\(6) & ( !\R.curInst\(5) & ( (!\R.curInst\(3) & ((!\R.curInst\(2)) # (\R.curInst\(4)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000110010001100000000000000000010001100100011001101100011011000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(2),
	datab => \ALT_INV_R.curInst\(3),
	datac => \ALT_INV_R.curInst\(4),
	datae => \ALT_INV_R.curInst\(6),
	dataf => \ALT_INV_R.curInst\(5),
	combout => \Mux34~0_combout\);

-- Location: IOIBUF_X80_Y0_N18
\avm_i_readdata[22]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(22),
	o => \avm_i_readdata[22]~input_o\);

-- Location: DDIOINCELL_X80_Y0_N31
\R.curInst[14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[22]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(14));

-- Location: IOIBUF_X80_Y0_N52
\avm_i_readdata[21]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(21),
	o => \avm_i_readdata[21]~input_o\);

-- Location: DDIOINCELL_X80_Y0_N65
\R.curInst[13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[21]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(13));

-- Location: IOIBUF_X78_Y0_N18
\avm_i_readdata[20]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(20),
	o => \avm_i_readdata[20]~input_o\);

-- Location: DDIOINCELL_X78_Y0_N31
\R.curInst[12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[20]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(12));

-- Location: LABCELL_X79_Y4_N0
\Mux0~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux0~0_combout\ = ( !\R.curInst\(12) & ( (!\R.curInst\(14) & !\R.curInst\(13)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1100000011000000110000001100000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.curInst\(14),
	datac => \ALT_INV_R.curInst\(13),
	dataf => \ALT_INV_R.curInst\(12),
	combout => \Mux0~0_combout\);

-- Location: LABCELL_X80_Y2_N42
\Mux11~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux11~0_combout\ = ( \R.curInst\(5) & ( \Mux0~0_combout\ & ( (!\R.curInst\(3) & (!\R.curInst\(2) & (\R.curInst\(4) & \R.curInst\(6)))) ) ) ) # ( !\R.curInst\(5) & ( \Mux0~0_combout\ & ( (\R.curInst\(3) & (\R.curInst\(2) & (!\R.curInst\(4) & 
-- !\R.curInst\(6)))) ) ) ) # ( !\R.curInst\(5) & ( !\Mux0~0_combout\ & ( (\R.curInst\(3) & (\R.curInst\(2) & (!\R.curInst\(4) & !\R.curInst\(6)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000000000000000000000000000000010000000000000000000000001000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(3),
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_R.curInst\(4),
	datad => \ALT_INV_R.curInst\(6),
	datae => \ALT_INV_R.curInst\(5),
	dataf => \ALT_INV_Mux0~0_combout\,
	combout => \Mux11~0_combout\);

-- Location: MLABCELL_X82_Y1_N39
\NxR~12\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR~12_combout\ = ( \R.ctrlState.Calc~q\ & ( \Mux11~0_combout\ & ( (!\Equal4~1_combout\) # ((!\R.ctrlState.ReadReg~q\ & !\Mux34~0_combout\)) ) ) ) # ( !\R.ctrlState.Calc~q\ & ( \Mux11~0_combout\ & ( (!\Equal4~1_combout\ & \R.ctrlState.ReadReg~q\) ) ) ) # 
-- ( \R.ctrlState.Calc~q\ & ( !\Mux11~0_combout\ & ( (!\Equal4~1_combout\) # ((!\Mux34~0_combout\) # (\R.ctrlState.ReadReg~q\)) ) ) ) # ( !\R.ctrlState.Calc~q\ & ( !\Mux11~0_combout\ & ( \R.ctrlState.ReadReg~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111111111111100111100001100000011001111110011001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Equal4~1_combout\,
	datac => \ALT_INV_R.ctrlState.ReadReg~q\,
	datad => \ALT_INV_Mux34~0_combout\,
	datae => \ALT_INV_R.ctrlState.Calc~q\,
	dataf => \ALT_INV_Mux11~0_combout\,
	combout => \NxR~12_combout\);

-- Location: FF_X82_Y1_N40
\R.ctrlState.Calc\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR~12_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.ctrlState.Calc~q\);

-- Location: LABCELL_X77_Y1_N15
\Mux53~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux53~0_combout\ = ( !\R.curInst\(2) & ( !\R.curInst\(3) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111000011110000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.curInst\(3),
	dataf => \ALT_INV_R.curInst\(2),
	combout => \Mux53~0_combout\);

-- Location: FF_X80_Y1_N40
\R.ctrlState.DataAccess0~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR~13_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.ctrlState.DataAccess0~DUPLICATE_q\);

-- Location: MLABCELL_X78_Y1_N45
\Mux50~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux50~0_combout\ = ( \R.curInst\(0) & ( (!\R.curInst\(6) & (!\R.curInst\(4))) # (\R.curInst\(6) & (\R.curInst\(4) & \R.curInst\(5))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000010001001100010011000100110001001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(6),
	datab => \ALT_INV_R.curInst\(4),
	datac => \ALT_INV_R.curInst\(5),
	dataf => \ALT_INV_R.curInst\(0),
	combout => \Mux50~0_combout\);

-- Location: LABCELL_X80_Y1_N39
\NxR~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR~13_combout\ = ( \Mux50~0_combout\ & ( (!\R.ctrlState.Calc~q\ & (\R.ctrlState.DataAccess0~DUPLICATE_q\ & ((!\Mux53~0_combout\) # (!\R.curInst\(1))))) # (\R.ctrlState.Calc~q\ & (\Mux53~0_combout\ & ((\R.curInst\(1))))) ) ) # ( !\Mux50~0_combout\ & ( 
-- (\R.ctrlState.DataAccess0~DUPLICATE_q\ & !\R.ctrlState.Calc~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100000000001100110000000000110010000001010011001000000101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux53~0_combout\,
	datab => \ALT_INV_R.ctrlState.DataAccess0~DUPLICATE_q\,
	datac => \ALT_INV_R.curInst\(1),
	datad => \ALT_INV_R.ctrlState.Calc~q\,
	dataf => \ALT_INV_Mux50~0_combout\,
	combout => \NxR~13_combout\);

-- Location: FF_X80_Y1_N41
\R.ctrlState.DataAccess0\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR~13_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.ctrlState.DataAccess0~q\);

-- Location: LABCELL_X77_Y5_N15
\Mux18~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux18~0_combout\ = ( \R.curInst\(5) & ( !\R.curInst\(4) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011110000111100001111000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.curInst\(4),
	dataf => \ALT_INV_R.curInst\(5),
	combout => \Mux18~0_combout\);

-- Location: LABCELL_X80_Y1_N6
\Mux53~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux53~1_combout\ = ( \Equal4~1_combout\ & ( \Mux53~0_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Mux53~0_combout\,
	dataf => \ALT_INV_Equal4~1_combout\,
	combout => \Mux53~1_combout\);

-- Location: LABCELL_X80_Y1_N27
\Mux53~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux53~2_combout\ = (\R.curInst\(4) & (\Mux53~1_combout\ & (\R.curInst\(5) & \R.curInst\(6))))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000001000000000000000100000000000000010000000000000001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(4),
	datab => \ALT_INV_Mux53~1_combout\,
	datac => \ALT_INV_R.curInst\(5),
	datad => \ALT_INV_R.curInst\(6),
	combout => \Mux53~2_combout\);

-- Location: IOIBUF_X80_Y0_N35
\avm_i_readdata[3]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(3),
	o => \avm_i_readdata[3]~input_o\);

-- Location: DDIOINCELL_X80_Y0_N48
\R.curInst[27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[3]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(27));

-- Location: IOIBUF_X80_Y0_N1
\avm_i_readdata[5]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(5),
	o => \avm_i_readdata[5]~input_o\);

-- Location: DDIOINCELL_X80_Y0_N14
\R.curInst[29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[5]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(29));

-- Location: IOIBUF_X74_Y0_N75
\avm_i_readdata[6]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(6),
	o => \avm_i_readdata[6]~input_o\);

-- Location: DDIOINCELL_X74_Y0_N88
\R.curInst[30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[6]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(30));

-- Location: IOIBUF_X74_Y0_N92
\avm_i_readdata[4]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(4),
	o => \avm_i_readdata[4]~input_o\);

-- Location: DDIOINCELL_X74_Y0_N105
\R.curInst[28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[4]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(28));

-- Location: IOIBUF_X74_Y0_N58
\avm_i_readdata[7]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(7),
	o => \avm_i_readdata[7]~input_o\);

-- Location: DDIOINCELL_X74_Y0_N71
\R.curInst[31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[7]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(31));

-- Location: LABCELL_X77_Y1_N12
\Equal2~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Equal2~0_combout\ = ( !\R.curInst\(31) & ( (!\R.curInst\(27) & (\R.curInst\(29) & (!\R.curInst\(30) & \R.curInst\(28)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000100000000000000010000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(27),
	datab => \ALT_INV_R.curInst\(29),
	datac => \ALT_INV_R.curInst\(30),
	datad => \ALT_INV_R.curInst\(28),
	dataf => \ALT_INV_R.curInst\(31),
	combout => \Equal2~0_combout\);

-- Location: IOIBUF_X82_Y0_N92
\avm_i_readdata[2]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(2),
	o => \avm_i_readdata[2]~input_o\);

-- Location: DDIOINCELL_X82_Y0_N105
\R.curInst[26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[2]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(26));

-- Location: IOIBUF_X66_Y0_N92
\avm_i_readdata[14]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(14),
	o => \avm_i_readdata[14]~input_o\);

-- Location: DDIOINCELL_X66_Y0_N105
\R.curInst[22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[14]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(22));

-- Location: IOIBUF_X70_Y0_N52
\avm_i_readdata[15]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(15),
	o => \avm_i_readdata[15]~input_o\);

-- Location: DDIOINCELL_X70_Y0_N65
\R.curInst[23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[15]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(23));

-- Location: IOIBUF_X74_Y0_N41
\avm_i_readdata[1]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(1),
	o => \avm_i_readdata[1]~input_o\);

-- Location: DDIOINCELL_X74_Y0_N54
\R.curInst[25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[1]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(25));

-- Location: IOIBUF_X72_Y0_N1
\avm_i_readdata[0]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(0),
	o => \avm_i_readdata[0]~input_o\);

-- Location: DDIOINCELL_X72_Y0_N14
\R.curInst[24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[0]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(24));

-- Location: LABCELL_X77_Y1_N36
\Equal2~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Equal2~1_combout\ = ( !\R.curInst\(25) & ( !\R.curInst\(24) & ( (!\R.curInst\(22) & !\R.curInst\(23)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010000010100000000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_R.curInst\(23),
	datae => \ALT_INV_R.curInst\(25),
	dataf => \ALT_INV_R.curInst\(24),
	combout => \Equal2~1_combout\);

-- Location: IOIBUF_X66_Y0_N58
\avm_i_readdata[13]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(13),
	o => \avm_i_readdata[13]~input_o\);

-- Location: DDIOINCELL_X66_Y0_N71
\R.curInst[21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[13]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(21));

-- Location: LABCELL_X77_Y1_N24
\Equal2~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Equal2~2_combout\ = ( \Equal2~1_combout\ & ( \R.curInst\(21) & ( ((!\Equal2~0_combout\) # (\R.curInst\(26))) # (\R.curInst\(20)) ) ) ) # ( !\Equal2~1_combout\ & ( \R.curInst\(21) ) ) # ( \Equal2~1_combout\ & ( !\R.curInst\(21) ) ) # ( !\Equal2~1_combout\ 
-- & ( !\R.curInst\(21) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111111111111111111111111111111111111101111111011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(20),
	datab => \ALT_INV_Equal2~0_combout\,
	datac => \ALT_INV_R.curInst\(26),
	datae => \ALT_INV_Equal2~1_combout\,
	dataf => \ALT_INV_R.curInst\(21),
	combout => \Equal2~2_combout\);

-- Location: LABCELL_X80_Y1_N0
\NxR~20\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR~20_combout\ = ( !\R.ctrlState.ReadReg~q\ & ( (!\R.ctrlState.Calc~q\ & (((\Equal2~2_combout\ & (!\R.ctrlState.DataAccess0~q\ & \R.ctrlState.Trap~q\))))) ) ) # ( \R.ctrlState.ReadReg~q\ & ( ((\Mux0~0_combout\ & (\Mux53~2_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000000000000000110000001100001010000000000000001100000011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.ctrlState.Calc~q\,
	datab => \ALT_INV_Mux0~0_combout\,
	datac => \ALT_INV_Mux53~2_combout\,
	datad => \ALT_INV_R.ctrlState.DataAccess0~q\,
	datae => \ALT_INV_R.ctrlState.ReadReg~q\,
	dataf => \ALT_INV_R.ctrlState.Trap~q\,
	datag => \ALT_INV_Equal2~2_combout\,
	combout => \NxR~20_combout\);

-- Location: FF_X80_Y1_N1
\R.ctrlState.Trap\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR~20_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.ctrlState.Trap~q\);

-- Location: LABCELL_X80_Y1_N30
\NxR~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR~18_combout\ = ( \Mux53~1_combout\ & ( (!\R.curInst\(4) & (\R.ctrlState.Calc~q\ & (\R.curInst\(6) & \R.curInst\(5)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000100000000000000010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(4),
	datab => \ALT_INV_R.ctrlState.Calc~q\,
	datac => \ALT_INV_R.curInst\(6),
	datad => \ALT_INV_R.curInst\(5),
	dataf => \ALT_INV_Mux53~1_combout\,
	combout => \NxR~18_combout\);

-- Location: FF_X80_Y1_N31
\R.ctrlState.CheckJump\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR~18_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.ctrlState.CheckJump~q\);

-- Location: LABCELL_X77_Y5_N12
\Mux154~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux154~0_combout\ = ( !\R.curInst\(5) & ( !\R.curInst\(6) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111100000000111111110000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \ALT_INV_R.curInst\(6),
	dataf => \ALT_INV_R.curInst\(5),
	combout => \Mux154~0_combout\);

-- Location: MLABCELL_X78_Y1_N15
\NxR~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR~4_combout\ = ( \Equal4~1_combout\ & ( \Mux154~0_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000111111110000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \ALT_INV_Mux154~0_combout\,
	dataf => \ALT_INV_Equal4~1_combout\,
	combout => \NxR~4_combout\);

-- Location: MLABCELL_X78_Y1_N18
\Mux12~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux12~0_combout\ = ( \NxR~4_combout\ & ( (!\R.curInst\(4) & (\R.curInst\(3) & \R.curInst\(2))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000011000000000000001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.curInst\(4),
	datac => \ALT_INV_R.curInst\(3),
	datad => \ALT_INV_R.curInst\(2),
	dataf => \ALT_INV_NxR~4_combout\,
	combout => \Mux12~0_combout\);

-- Location: MLABCELL_X78_Y1_N0
\NxR~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR~14_combout\ = ( \R.ctrlState.CheckJump~q\ & ( \Mux12~0_combout\ & ( ((!\R.ctrlState.DataAccess0~DUPLICATE_q\ & !\R.ctrlState.Calc~q\)) # (\R.ctrlState.ReadReg~q\) ) ) ) # ( !\R.ctrlState.CheckJump~q\ & ( \Mux12~0_combout\ & ( \R.ctrlState.ReadReg~q\ 
-- ) ) ) # ( \R.ctrlState.CheckJump~q\ & ( !\Mux12~0_combout\ & ( (!\R.ctrlState.DataAccess0~DUPLICATE_q\ & (!\R.ctrlState.ReadReg~q\ & !\R.ctrlState.Calc~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110000000000000000001111000011111100111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.ctrlState.DataAccess0~DUPLICATE_q\,
	datac => \ALT_INV_R.ctrlState.ReadReg~q\,
	datad => \ALT_INV_R.ctrlState.Calc~q\,
	datae => \ALT_INV_R.ctrlState.CheckJump~q\,
	dataf => \ALT_INV_Mux12~0_combout\,
	combout => \NxR~14_combout\);

-- Location: FF_X78_Y1_N2
\R.ctrlState.Wait0\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR~14_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.ctrlState.Wait0~q\);

-- Location: LABCELL_X77_Y1_N21
\NxR~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR~0_combout\ = ( \Equal2~2_combout\ & ( !\R.ctrlState.Wait0~q\ ) ) # ( !\Equal2~2_combout\ & ( (!\R.ctrlState.Trap~q\ & !\R.ctrlState.Wait0~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111000000000000111100000000000011111111000000001111111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.ctrlState.Trap~q\,
	datad => \ALT_INV_R.ctrlState.Wait0~q\,
	dataf => \ALT_INV_Equal2~2_combout\,
	combout => \NxR~0_combout\);

-- Location: MLABCELL_X78_Y1_N54
\NxR~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR~1_combout\ = ( \NxR~0_combout\ & ( \Mux53~1_combout\ & ( (!\Mux18~0_combout\) # ((!\R.ctrlState.DataAccess0~DUPLICATE_q\) # ((\R.ctrlState.Calc~q\) # (\R.curInst\(6)))) ) ) ) # ( !\NxR~0_combout\ & ( \Mux53~1_combout\ & ( 
-- ((\R.ctrlState.DataAccess0~DUPLICATE_q\ & ((!\Mux18~0_combout\) # (\R.curInst\(6))))) # (\R.ctrlState.Calc~q\) ) ) ) # ( \NxR~0_combout\ & ( !\Mux53~1_combout\ ) ) # ( !\NxR~0_combout\ & ( !\Mux53~1_combout\ & ( (\R.ctrlState.Calc~q\) # 
-- (\R.ctrlState.DataAccess0~DUPLICATE_q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001111111111111111111111111100100011111111111110111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux18~0_combout\,
	datab => \ALT_INV_R.ctrlState.DataAccess0~DUPLICATE_q\,
	datac => \ALT_INV_R.curInst\(6),
	datad => \ALT_INV_R.ctrlState.Calc~q\,
	datae => \ALT_INV_NxR~0_combout\,
	dataf => \ALT_INV_Mux53~1_combout\,
	combout => \NxR~1_combout\);

-- Location: FF_X78_Y1_N55
\R.ctrlState.Wait1\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR~1_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.ctrlState.Wait1~q\);

-- Location: LABCELL_X75_Y3_N0
\vAluSrc1~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluSrc1~0_combout\ = ( !\R.curInst\(3) & ( (!\R.curInst\(6) & \R.curInst\(4)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011001100000000001100110000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.curInst\(6),
	datad => \ALT_INV_R.curInst\(4),
	dataf => \ALT_INV_R.curInst\(3),
	combout => \vAluSrc1~0_combout\);

-- Location: LABCELL_X77_Y5_N9
\Mux123~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux123~0_combout\ = ( \R.curInst\(5) & ( (\R.curInst\(2) & \R.curInst\(6)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000010101010000000001010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(2),
	datad => \ALT_INV_R.curInst\(6),
	dataf => \ALT_INV_R.curInst\(5),
	combout => \Mux123~0_combout\);

-- Location: LABCELL_X80_Y1_N33
\NxR~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR~2_combout\ = ( \Mux123~0_combout\ & ( (\R.ctrlState.Calc~q\ & (\Equal4~1_combout\ & ((!\R.curInst\(4)) # (\vAluSrc1~0_combout\)))) ) ) # ( !\Mux123~0_combout\ & ( (\R.ctrlState.Calc~q\ & (\Equal4~1_combout\ & \vAluSrc1~0_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000011000000000000001100000010000000110000001000000011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(4),
	datab => \ALT_INV_R.ctrlState.Calc~q\,
	datac => \ALT_INV_Equal4~1_combout\,
	datad => \ALT_INV_vAluSrc1~0_combout\,
	dataf => \ALT_INV_Mux123~0_combout\,
	combout => \NxR~2_combout\);

-- Location: LABCELL_X80_Y1_N36
\NxR~15\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR~15_combout\ = ( \NxR~4_combout\ & ( (\Mux53~0_combout\ & (\R.ctrlState.DataAccess0~DUPLICATE_q\ & !\R.curInst\(4))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000010000000100000001000000010000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux53~0_combout\,
	datab => \ALT_INV_R.ctrlState.DataAccess0~DUPLICATE_q\,
	datac => \ALT_INV_R.curInst\(4),
	dataf => \ALT_INV_NxR~4_combout\,
	combout => \NxR~15_combout\);

-- Location: LABCELL_X80_Y1_N15
\NxR~16\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR~16_combout\ = (!\R.ctrlState.Calc~q\ & \NxR~15_combout\)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011110000000000001111000000000000111100000000000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.ctrlState.Calc~q\,
	datad => \ALT_INV_NxR~15_combout\,
	combout => \NxR~16_combout\);

-- Location: FF_X80_Y1_N16
\R.ctrlState.DataAccess1\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR~16_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.ctrlState.DataAccess1~q\);

-- Location: LABCELL_X80_Y1_N9
\NxR~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR~3_combout\ = ( \R.ctrlState.DataAccess1~q\ & ( ((!\R.ctrlState.Calc~q\ & ((!\R.ctrlState.DataAccess0~q\) # (\Mux53~2_combout\)))) # (\NxR~2_combout\) ) ) # ( !\R.ctrlState.DataAccess1~q\ & ( ((!\R.ctrlState.Calc~q\ & (\R.ctrlState.DataAccess0~q\ & 
-- \Mux53~2_combout\))) # (\NxR~2_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101011101010101010101110111010101110111011101010111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_NxR~2_combout\,
	datab => \ALT_INV_R.ctrlState.Calc~q\,
	datac => \ALT_INV_R.ctrlState.DataAccess0~q\,
	datad => \ALT_INV_Mux53~2_combout\,
	dataf => \ALT_INV_R.ctrlState.DataAccess1~q\,
	combout => \NxR~3_combout\);

-- Location: FF_X80_Y1_N11
\R.ctrlState.WriteReg\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR~3_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.ctrlState.WriteReg~q\);

-- Location: LABCELL_X80_Y1_N45
\Comb~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb~0_combout\ = ( \R.ctrlState.WriteReg~q\ ) # ( !\R.ctrlState.WriteReg~q\ & ( !\R.ctrlState.Wait1~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111000011110000111100001111000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.ctrlState.Wait1~q\,
	dataf => \ALT_INV_R.ctrlState.WriteReg~q\,
	combout => \Comb~0_combout\);

-- Location: LABCELL_X80_Y1_N57
\NxR~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR~17_combout\ = (!\R.ctrlState.Calc~q\ & (!\R.ctrlState.DataAccess0~q\ & \Comb~0_combout\))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011000000000000001100000000000000110000000000000011000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.ctrlState.Calc~q\,
	datac => \ALT_INV_R.ctrlState.DataAccess0~q\,
	datad => \ALT_INV_Comb~0_combout\,
	combout => \NxR~17_combout\);

-- Location: FF_X80_Y1_N59
\R.ctrlState.Fetch\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR~17_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.ctrlState.Fetch~q\);

-- Location: FF_X74_Y4_N35
\R.ctrlState.ReadReg\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.ctrlState.Fetch~q\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.ctrlState.ReadReg~q\);

-- Location: LABCELL_X74_Y4_N36
\vAluSrc2~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluSrc2~0_combout\ = ( \R.curInst\(1) & ( (\R.curInst\(0) & \R.ctrlState.ReadReg~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000011000000110000001100000011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.curInst\(0),
	datac => \ALT_INV_R.ctrlState.ReadReg~q\,
	dataf => \ALT_INV_R.curInst\(1),
	combout => \vAluSrc2~0_combout\);

-- Location: LABCELL_X74_Y4_N30
\vAluSrc2~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluSrc2~1_combout\ = ( \vAluSrc2~0_combout\ & ( \R.curInst\(6) & ( (!\R.curInst\(4) & (\R.curInst\(2) & (\R.curInst\(5) & !\R.curInst\(3)))) ) ) ) # ( \vAluSrc2~0_combout\ & ( !\R.curInst\(6) & ( (!\R.curInst\(3) & ((!\R.curInst\(4) & (!\R.curInst\(2))) 
-- # (\R.curInst\(4) & ((!\R.curInst\(5)) # (\R.curInst\(2)))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110110010000000000000000000000000000001000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(4),
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_R.curInst\(5),
	datad => \ALT_INV_R.curInst\(3),
	datae => \ALT_INV_vAluSrc2~0_combout\,
	dataf => \ALT_INV_R.curInst\(6),
	combout => \vAluSrc2~1_combout\);

-- Location: LABCELL_X81_Y1_N42
\~GND\ : cyclonev_lcell_comb
-- Equation(s):
-- \~GND~combout\ = GND

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	combout => \~GND~combout\);

-- Location: FF_X80_Y1_N38
\R.memToReg\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR~15_combout\,
	asdata => \~GND~combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sclr => \R.ctrlState.Fetch~q\,
	sload => \R.ctrlState.ReadReg~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.memToReg~q\);

-- Location: IOIBUF_X70_Y0_N35
\avm_d_readdata[24]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(24),
	o => \avm_d_readdata[24]~input_o\);

-- Location: LABCELL_X81_Y1_N39
\Comb:vRegWriteData[0]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[0]~0_combout\ = ( !\R.curInst\(12) & ( \R.curInst\(13) & ( (\R.memToReg~q\ & (\avm_d_readdata[24]~input_o\ & !\R.curInst\(14))) ) ) ) # ( \R.curInst\(12) & ( !\R.curInst\(13) & ( (\R.memToReg~q\ & \avm_d_readdata[24]~input_o\) ) ) ) # 
-- ( !\R.curInst\(12) & ( !\R.curInst\(13) & ( (\R.memToReg~q\ & \avm_d_readdata[24]~input_o\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100010001000100010001000100010000000100000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.memToReg~q\,
	datab => \ALT_INV_avm_d_readdata[24]~input_o\,
	datac => \ALT_INV_R.curInst\(14),
	datae => \ALT_INV_R.curInst\(12),
	dataf => \ALT_INV_R.curInst\(13),
	combout => \Comb:vRegWriteData[0]~0_combout\);

-- Location: LABCELL_X79_Y4_N39
\NxR~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR~5_combout\ = ( !\Mux12~0_combout\ & ( \R.ctrlState.ReadReg~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101010101010101010100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.ctrlState.ReadReg~q\,
	dataf => \ALT_INV_Mux12~0_combout\,
	combout => \NxR~5_combout\);

-- Location: FF_X79_Y4_N41
\R.aluCalc\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR~5_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sclr => \R.ctrlState.Fetch~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluCalc~q\);

-- Location: LABCELL_X75_Y4_N3
\Mux124~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux124~0_combout\ = ( \R.curInst\(31) & ( (!\R.curInst\(5) & !\R.curInst\(2)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000010001000100010001000100010001000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(5),
	datab => \ALT_INV_R.curInst\(2),
	dataf => \ALT_INV_R.curInst\(31),
	combout => \Mux124~0_combout\);

-- Location: LABCELL_X74_Y4_N48
\Mux123~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux123~1_combout\ = ( \R.curInst\(2) & ( \R.curInst\(31) & ( (!\R.curInst\(4) & (\R.curInst\(6) & \R.curInst\(5))) ) ) ) # ( !\R.curInst\(2) & ( \R.curInst\(31) & ( (!\R.curInst\(4) & (!\R.curInst\(3) & ((!\R.curInst\(6)) # (\R.curInst\(5))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000010001010000000000000001000000010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(4),
	datab => \ALT_INV_R.curInst\(6),
	datac => \ALT_INV_R.curInst\(5),
	datad => \ALT_INV_R.curInst\(3),
	datae => \ALT_INV_R.curInst\(2),
	dataf => \ALT_INV_R.curInst\(31),
	combout => \Mux123~1_combout\);

-- Location: LABCELL_X75_Y4_N21
\Mux131~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux131~0_combout\ = ( \vAluSrc1~0_combout\ & ( (((\R.curInst\(2) & \R.curInst\(23))) # (\Mux123~1_combout\)) # (\Mux124~0_combout\) ) ) # ( !\vAluSrc1~0_combout\ & ( \Mux123~1_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111000000001111111101010111111111110101011111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux124~0_combout\,
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_R.curInst\(23),
	datad => \ALT_INV_Mux123~1_combout\,
	dataf => \ALT_INV_vAluSrc1~0_combout\,
	combout => \Mux131~0_combout\);

-- Location: MLABCELL_X78_Y1_N51
\Comb~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb~1_combout\ = ( \Equal4~1_combout\ & ( (\vAluSrc1~0_combout\ & (\R.curInst\(30) & (\R.curInst\(5) & !\R.curInst\(2)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000001000000000000000100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluSrc1~0_combout\,
	datab => \ALT_INV_R.curInst\(30),
	datac => \ALT_INV_R.curInst\(5),
	datad => \ALT_INV_R.curInst\(2),
	dataf => \ALT_INV_Equal4~1_combout\,
	combout => \Comb~1_combout\);

-- Location: LABCELL_X77_Y1_N0
\Mux18~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux18~1_combout\ = ( \R.curInst\(5) & ( \Comb~1_combout\ & ( (!\R.curInst\(4) & (\R.aluOp.ALUOpSub~q\ & ((\R.curInst\(2))))) # (\R.curInst\(4) & (((\Mux0~0_combout\ & !\R.curInst\(2))))) ) ) ) # ( !\R.curInst\(5) & ( \Comb~1_combout\ & ( 
-- (\R.aluOp.ALUOpSub~q\ & (!\R.curInst\(4) & \R.curInst\(2))) ) ) ) # ( \R.curInst\(5) & ( !\Comb~1_combout\ & ( (\R.aluOp.ALUOpSub~q\ & (!\R.curInst\(4) & \R.curInst\(2))) ) ) ) # ( !\R.curInst\(5) & ( !\Comb~1_combout\ & ( (\R.aluOp.ALUOpSub~q\ & 
-- (!\R.curInst\(4) & \R.curInst\(2))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001000100000000000100010000000000010001000000001101000100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datab => \ALT_INV_R.curInst\(4),
	datac => \ALT_INV_Mux0~0_combout\,
	datad => \ALT_INV_R.curInst\(2),
	datae => \ALT_INV_R.curInst\(5),
	dataf => \ALT_INV_Comb~1_combout\,
	combout => \Mux18~1_combout\);

-- Location: MLABCELL_X78_Y1_N30
\Mux18~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux18~2_combout\ = ( \R.aluOp.ALUOpSub~q\ & ( \Mux18~1_combout\ & ( (!\R.curInst\(6)) # ((!\R.curInst\(2)) # (!\Mux18~0_combout\)) ) ) ) # ( !\R.aluOp.ALUOpSub~q\ & ( \Mux18~1_combout\ & ( (!\R.curInst\(3) & ((!\R.curInst\(6)) # ((!\R.curInst\(2) & 
-- \Mux18~0_combout\)))) ) ) ) # ( \R.aluOp.ALUOpSub~q\ & ( !\Mux18~1_combout\ & ( (!\R.curInst\(6) & (((\R.curInst\(3))))) # (\R.curInst\(6) & ((!\R.curInst\(2)) # ((!\Mux18~0_combout\)))) ) ) ) # ( !\R.aluOp.ALUOpSub~q\ & ( !\Mux18~1_combout\ & ( 
-- (\R.curInst\(6) & (!\R.curInst\(2) & (\Mux18~0_combout\ & !\R.curInst\(3)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010000000000010101001111111010101110000000001111111011111110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(6),
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_Mux18~0_combout\,
	datad => \ALT_INV_R.curInst\(3),
	datae => \ALT_INV_R.aluOp.ALUOpSub~q\,
	dataf => \ALT_INV_Mux18~1_combout\,
	combout => \Mux18~2_combout\);

-- Location: FF_X78_Y1_N31
\R.aluOp.ALUOpSub\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Mux18~2_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \vAluSrc2~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluOp.ALUOpSub~q\);

-- Location: MLABCELL_X78_Y1_N27
\Mux17~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux17~0_combout\ = ( \R.aluOp.ALUOpAdd~q\ & ( (\R.curInst\(4) & (!\R.curInst\(2) & ((!\Mux0~0_combout\) # (\Comb~1_combout\)))) ) ) # ( !\R.aluOp.ALUOpAdd~q\ & ( (!\R.curInst\(4) & (((\R.curInst\(2))))) # (\R.curInst\(4) & (!\R.curInst\(2) & 
-- ((!\Mux0~0_combout\) # (\Comb~1_combout\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011110000011100001111000001110000110000000100000011000000010000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Comb~1_combout\,
	datab => \ALT_INV_R.curInst\(4),
	datac => \ALT_INV_R.curInst\(2),
	datad => \ALT_INV_Mux0~0_combout\,
	dataf => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	combout => \Mux17~0_combout\);

-- Location: MLABCELL_X78_Y1_N6
\Mux17~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux17~1_combout\ = ( \Mux17~0_combout\ & ( \R.aluOp.ALUOpAdd~q\ & ( (!\R.curInst\(6) & (((\R.curInst\(3))))) # (\R.curInst\(6) & ((!\Mux18~0_combout\) # (!\R.curInst\(2) $ (!\R.curInst\(3))))) ) ) ) # ( !\Mux17~0_combout\ & ( \R.aluOp.ALUOpAdd~q\ & ( 
-- (!\R.curInst\(6)) # ((!\Mux18~0_combout\) # (!\R.curInst\(2) $ (!\R.curInst\(3)))) ) ) ) # ( \Mux17~0_combout\ & ( !\R.aluOp.ALUOpAdd~q\ & ( (\R.curInst\(6) & (\R.curInst\(2) & (\Mux18~0_combout\ & !\R.curInst\(3)))) ) ) ) # ( !\Mux17~0_combout\ & ( 
-- !\R.aluOp.ALUOpAdd~q\ & ( (!\R.curInst\(3) & ((!\R.curInst\(6)) # ((\R.curInst\(2) & \Mux18~0_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010101100000000000000010000000011111011111111100101000111111110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(6),
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_Mux18~0_combout\,
	datad => \ALT_INV_R.curInst\(3),
	datae => \ALT_INV_Mux17~0_combout\,
	dataf => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	combout => \Mux17~1_combout\);

-- Location: MLABCELL_X78_Y1_N48
\R.aluOp.ALUOpAdd_NEW364\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.aluOp.ALUOpAdd_OTERM365\ = ( \Mux17~1_combout\ & ( (\R.aluOp.ALUOpAdd~q\) # (\vAluSrc2~0_combout\) ) ) # ( !\Mux17~1_combout\ & ( (!\vAluSrc2~0_combout\ & \R.aluOp.ALUOpAdd~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011110000000000001111000000001111111111110000111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_vAluSrc2~0_combout\,
	datad => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	dataf => \ALT_INV_Mux17~1_combout\,
	combout => \R.aluOp.ALUOpAdd_OTERM365\);

-- Location: FF_X78_Y1_N50
\R.aluOp.ALUOpAdd\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \R.aluOp.ALUOpAdd_OTERM365\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluOp.ALUOpAdd~q\);

-- Location: LABCELL_X74_Y4_N39
\vAluSrc1~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluSrc1~2_combout\ = ( !\R.curInst\(5) & ( (\vAluSrc1~0_combout\ & (\R.curInst\(2) & \vAluSrc2~0_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000101000000000000010100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluSrc1~0_combout\,
	datac => \ALT_INV_R.curInst\(2),
	datad => \ALT_INV_vAluSrc2~0_combout\,
	dataf => \ALT_INV_R.curInst\(5),
	combout => \vAluSrc1~2_combout\);

-- Location: LABCELL_X74_Y4_N18
\vAluSrc1~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluSrc1~1_combout\ = ( \R.curInst\(5) & ( (\vAluSrc1~0_combout\ & (\R.curInst\(2) & \vAluSrc2~0_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000100010000000000010001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluSrc1~0_combout\,
	datab => \ALT_INV_R.curInst\(2),
	datad => \ALT_INV_vAluSrc2~0_combout\,
	dataf => \ALT_INV_R.curInst\(5),
	combout => \vAluSrc1~1_combout\);

-- Location: IOIBUF_X64_Y0_N35
\avm_i_readdata[10]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(10),
	o => \avm_i_readdata[10]~input_o\);

-- Location: DDIOINCELL_X64_Y0_N48
\R.curInst[18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[10]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(18));

-- Location: IOIBUF_X66_Y0_N41
\avm_i_readdata[11]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(11),
	o => \avm_i_readdata[11]~input_o\);

-- Location: DDIOINCELL_X66_Y0_N54
\R.curInst[19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[11]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(19));

-- Location: IOIBUF_X68_Y0_N1
\avm_i_readdata[19]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(19),
	o => \avm_i_readdata[19]~input_o\);

-- Location: DDIOINCELL_X68_Y0_N14
\R.curInst[11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[19]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(11));

-- Location: IOIBUF_X68_Y0_N35
\avm_i_readdata[18]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(18),
	o => \avm_i_readdata[18]~input_o\);

-- Location: DDIOINCELL_X68_Y0_N48
\R.curInst[10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[18]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(10));

-- Location: IOIBUF_X68_Y0_N18
\avm_i_readdata[17]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(17),
	o => \avm_i_readdata[17]~input_o\);

-- Location: DDIOINCELL_X68_Y0_N31
\R.curInst[9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[17]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(9));

-- Location: IOIBUF_X68_Y0_N52
\avm_i_readdata[16]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(16),
	o => \avm_i_readdata[16]~input_o\);

-- Location: DDIOINCELL_X68_Y0_N65
\R.curInst[8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[16]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(8));

-- Location: LABCELL_X74_Y1_N54
\Mux31~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux31~0_combout\ = ( !\R.curInst\(9) & ( !\R.curInst\(8) & ( (!\R.curInst\(7) & (!\R.curInst\(11) & !\R.curInst\(10))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000000010000000000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(7),
	datab => \ALT_INV_R.curInst\(11),
	datac => \ALT_INV_R.curInst\(10),
	datae => \ALT_INV_R.curInst\(9),
	dataf => \ALT_INV_R.curInst\(8),
	combout => \Mux31~0_combout\);

-- Location: LABCELL_X80_Y1_N54
\NxR~19\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR~19_combout\ = ( \Mux31~0_combout\ & ( (\R.curInst\(13) & (\R.ctrlState.Calc~q\ & \Mux53~2_combout\)) ) ) # ( !\Mux31~0_combout\ & ( (\R.ctrlState.Calc~q\ & (\Mux53~2_combout\ & ((\R.curInst\(12)) # (\R.curInst\(13))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000010011000000000001001100000000000100010000000000010001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(13),
	datab => \ALT_INV_R.ctrlState.Calc~q\,
	datac => \ALT_INV_R.curInst\(12),
	datad => \ALT_INV_Mux53~2_combout\,
	dataf => \ALT_INV_Mux31~0_combout\,
	combout => \NxR~19_combout\);

-- Location: FF_X80_Y1_N56
\R.csrRead\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR~19_combout\,
	asdata => \~GND~combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sclr => \R.ctrlState.Fetch~q\,
	sload => \R.ctrlState.ReadReg~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.csrRead~q\);

-- Location: LABCELL_X80_Y1_N18
\R.regWriteEn~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.regWriteEn~1_combout\ = ( \Mux53~2_combout\ & ( !\NxR~2_combout\ & ( ((!\R.ctrlState.DataAccess0~DUPLICATE_q\ & ((!\R.ctrlState.DataAccess1~q\))) # (\R.ctrlState.DataAccess0~DUPLICATE_q\ & (!\R.csrRead~q\))) # (\R.ctrlState.Calc~q\) ) ) ) # ( 
-- !\Mux53~2_combout\ & ( !\NxR~2_combout\ & ( (!\R.ctrlState.DataAccess1~q\) # ((\R.ctrlState.Calc~q\) # (\R.ctrlState.DataAccess0~DUPLICATE_q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1100111111111111110010101111111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.csrRead~q\,
	datab => \ALT_INV_R.ctrlState.DataAccess1~q\,
	datac => \ALT_INV_R.ctrlState.DataAccess0~DUPLICATE_q\,
	datad => \ALT_INV_R.ctrlState.Calc~q\,
	datae => \ALT_INV_Mux53~2_combout\,
	dataf => \ALT_INV_NxR~2_combout\,
	combout => \R.regWriteEn~1_combout\);

-- Location: LABCELL_X80_Y1_N48
\R.regWriteEn~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.regWriteEn~0_combout\ = ( \Mux53~2_combout\ & ( \R.ctrlState.WriteReg~q\ & ( (!\R.ctrlState.ReadReg~q\ & (!\R.ctrlState.Calc~q\ & !\R.ctrlState.Fetch~q\)) ) ) ) # ( !\Mux53~2_combout\ & ( \R.ctrlState.WriteReg~q\ & ( (!\R.ctrlState.ReadReg~q\ & 
-- (!\R.ctrlState.Calc~q\ & (!\R.ctrlState.DataAccess0~DUPLICATE_q\ & !\R.ctrlState.Fetch~q\))) ) ) ) # ( \Mux53~2_combout\ & ( !\R.ctrlState.WriteReg~q\ & ( (!\R.ctrlState.ReadReg~q\ & (!\R.ctrlState.Calc~q\ & (\R.ctrlState.DataAccess0~DUPLICATE_q\ & 
-- !\R.ctrlState.Fetch~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000010000000000010000000000000001000100000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.ctrlState.ReadReg~q\,
	datab => \ALT_INV_R.ctrlState.Calc~q\,
	datac => \ALT_INV_R.ctrlState.DataAccess0~DUPLICATE_q\,
	datad => \ALT_INV_R.ctrlState.Fetch~q\,
	datae => \ALT_INV_Mux53~2_combout\,
	dataf => \ALT_INV_R.ctrlState.WriteReg~q\,
	combout => \R.regWriteEn~0_combout\);

-- Location: LABCELL_X80_Y1_N12
\R.regWriteEn~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.regWriteEn~2_combout\ = ( \R.regWriteEn~0_combout\ & ( (!\R.ctrlState.ReadReg~q\ & (!\R.ctrlState.Fetch~q\ & !\R.regWriteEn~1_combout\)) ) ) # ( !\R.regWriteEn~0_combout\ & ( ((!\R.ctrlState.ReadReg~q\ & (!\R.ctrlState.Fetch~q\ & 
-- !\R.regWriteEn~1_combout\))) # (\R.regWriteEn~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000000011111111100000001111111110000000100000001000000010000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.ctrlState.ReadReg~q\,
	datab => \ALT_INV_R.ctrlState.Fetch~q\,
	datac => \ALT_INV_R.regWriteEn~1_combout\,
	datad => \ALT_INV_R.regWriteEn~q\,
	dataf => \ALT_INV_R.regWriteEn~0_combout\,
	combout => \R.regWriteEn~2_combout\);

-- Location: FF_X80_Y1_N14
\R.regWriteEn\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \R.regWriteEn~2_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteEn~q\);

-- Location: LABCELL_X63_Y3_N51
\Decoder0~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~11_combout\ = ( \R.curInst\(9) & ( !\R.curInst\(8) & ( (\R.regWriteEn~q\ & (\R.curInst\(7) & (!\R.curInst\(10) & \R.curInst\(11)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000001000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.regWriteEn~q\,
	datab => \ALT_INV_R.curInst\(7),
	datac => \ALT_INV_R.curInst\(10),
	datad => \ALT_INV_R.curInst\(11),
	datae => \ALT_INV_R.curInst\(9),
	dataf => \ALT_INV_R.curInst\(8),
	combout => \Decoder0~11_combout\);

-- Location: FF_X64_Y1_N50
\RegFile[21][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(23),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][23]~q\);

-- Location: LABCELL_X71_Y3_N30
\Decoder0~12\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~12_combout\ = ( \R.curInst\(11) & ( \R.curInst\(8) & ( (!\R.curInst\(10) & (\R.curInst\(9) & (\R.regWriteEn~q\ & \R.curInst\(7)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000000000000000010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(10),
	datab => \ALT_INV_R.curInst\(9),
	datac => \ALT_INV_R.regWriteEn~q\,
	datad => \ALT_INV_R.curInst\(7),
	datae => \ALT_INV_R.curInst\(11),
	dataf => \ALT_INV_R.curInst\(8),
	combout => \Decoder0~12_combout\);

-- Location: FF_X70_Y3_N14
\RegFile[23][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(23),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][23]~q\);

-- Location: LABCELL_X71_Y1_N18
\RegFile[22][23]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[22][23]~feeder_combout\ = ( \R.regWriteData\(23) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(23),
	combout => \RegFile[22][23]~feeder_combout\);

-- Location: LABCELL_X68_Y5_N51
\Decoder0~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~14_combout\ = ( \R.curInst\(8) & ( \R.curInst\(11) & ( (!\R.curInst\(10) & (\R.curInst\(9) & (\R.regWriteEn~q\ & !\R.curInst\(7)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000000001000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(10),
	datab => \ALT_INV_R.curInst\(9),
	datac => \ALT_INV_R.regWriteEn~q\,
	datad => \ALT_INV_R.curInst\(7),
	datae => \ALT_INV_R.curInst\(8),
	dataf => \ALT_INV_R.curInst\(11),
	combout => \Decoder0~14_combout\);

-- Location: FF_X71_Y1_N19
\RegFile[22][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[22][23]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][23]~q\);

-- Location: IOIBUF_X64_Y0_N1
\avm_i_readdata[9]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(9),
	o => \avm_i_readdata[9]~input_o\);

-- Location: DDIOINCELL_X64_Y0_N14
\R.curInst[17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[9]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(17));

-- Location: IOIBUF_X64_Y0_N18
\avm_i_readdata[8]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(8),
	o => \avm_i_readdata[8]~input_o\);

-- Location: DDIOINCELL_X64_Y0_N31
\R.curInst[16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[8]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(16));

-- Location: LABCELL_X63_Y3_N18
\Decoder0~24\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~24_combout\ = ( \R.curInst\(7) & ( \R.curInst\(8) & ( (\R.regWriteEn~q\ & (!\R.curInst\(9) & (\R.curInst\(11) & !\R.curInst\(10)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000000010000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.regWriteEn~q\,
	datab => \ALT_INV_R.curInst\(9),
	datac => \ALT_INV_R.curInst\(11),
	datad => \ALT_INV_R.curInst\(10),
	datae => \ALT_INV_R.curInst\(7),
	dataf => \ALT_INV_R.curInst\(8),
	combout => \Decoder0~24_combout\);

-- Location: FF_X70_Y3_N50
\RegFile[19][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(23),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][23]~q\);

-- Location: LABCELL_X68_Y5_N27
\Decoder0~23\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~23_combout\ = ( \R.curInst\(11) & ( !\R.curInst\(10) & ( (!\R.curInst\(9) & (!\R.curInst\(8) & (\R.regWriteEn~q\ & \R.curInst\(7)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000100000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(9),
	datab => \ALT_INV_R.curInst\(8),
	datac => \ALT_INV_R.regWriteEn~q\,
	datad => \ALT_INV_R.curInst\(7),
	datae => \ALT_INV_R.curInst\(11),
	dataf => \ALT_INV_R.curInst\(10),
	combout => \Decoder0~23_combout\);

-- Location: FF_X64_Y1_N26
\RegFile[17][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(23),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][23]~q\);

-- Location: LABCELL_X63_Y3_N30
\Decoder0~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~26_combout\ = ( \R.curInst\(8) & ( !\R.curInst\(10) & ( (\R.regWriteEn~q\ & (!\R.curInst\(7) & (!\R.curInst\(9) & \R.curInst\(11)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000100000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.regWriteEn~q\,
	datab => \ALT_INV_R.curInst\(7),
	datac => \ALT_INV_R.curInst\(9),
	datad => \ALT_INV_R.curInst\(11),
	datae => \ALT_INV_R.curInst\(8),
	dataf => \ALT_INV_R.curInst\(10),
	combout => \Decoder0~26_combout\);

-- Location: FF_X59_Y3_N46
\RegFile[18][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(23),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][23]~q\);

-- Location: IOIBUF_X64_Y0_N52
\avm_i_readdata[23]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_readdata(23),
	o => \avm_i_readdata[23]~input_o\);

-- Location: DDIOINCELL_X64_Y0_N65
\R.curInst[15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \avm_i_readdata[23]~input_o\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curInst\(15));

-- Location: LABCELL_X64_Y1_N21
\RegFile[16][23]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[16][23]~feeder_combout\ = ( \R.regWriteData\(23) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(23),
	combout => \RegFile[16][23]~feeder_combout\);

-- Location: LABCELL_X68_Y5_N33
\Decoder0~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~25_combout\ = ( !\R.curInst\(8) & ( \R.curInst\(11) & ( (!\R.curInst\(10) & (!\R.curInst\(9) & (\R.regWriteEn~q\ & !\R.curInst\(7)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000001000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(10),
	datab => \ALT_INV_R.curInst\(9),
	datac => \ALT_INV_R.regWriteEn~q\,
	datad => \ALT_INV_R.curInst\(7),
	datae => \ALT_INV_R.curInst\(8),
	dataf => \ALT_INV_R.curInst\(11),
	combout => \Decoder0~25_combout\);

-- Location: FF_X64_Y1_N22
\RegFile[16][23]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[16][23]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][23]~DUPLICATE_q\);

-- Location: LABCELL_X70_Y3_N48
\Mux67~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux67~18_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[16][23]~DUPLICATE_q\))) # (\R.curInst\(15) & (\RegFile[17][23]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[18][23]~q\))) # (\R.curInst\(15) & (\RegFile[19][23]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[19][23]~q\,
	datab => \ALT_INV_RegFile[17][23]~q\,
	datac => \ALT_INV_RegFile[18][23]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][23]~DUPLICATE_q\,
	combout => \Mux67~18_combout\);

-- Location: LABCELL_X75_Y1_N21
\RegFile[20][23]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[20][23]~feeder_combout\ = ( \R.regWriteData\(23) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(23),
	combout => \RegFile[20][23]~feeder_combout\);

-- Location: LABCELL_X68_Y5_N18
\Decoder0~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~13_combout\ = ( !\R.curInst\(10) & ( !\R.curInst\(8) & ( (\R.curInst\(11) & (\R.curInst\(9) & (!\R.curInst\(7) & \R.regWriteEn~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000010000000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(11),
	datab => \ALT_INV_R.curInst\(9),
	datac => \ALT_INV_R.curInst\(7),
	datad => \ALT_INV_R.regWriteEn~q\,
	datae => \ALT_INV_R.curInst\(10),
	dataf => \ALT_INV_R.curInst\(8),
	combout => \Decoder0~13_combout\);

-- Location: FF_X75_Y1_N22
\RegFile[20][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[20][23]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][23]~q\);

-- Location: LABCELL_X70_Y3_N12
\Mux67~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux67~5_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux67~18_combout\)))) # (\R.curInst\(17) & ((!\Mux67~18_combout\ & ((\RegFile[20][23]~q\))) # (\Mux67~18_combout\ & (\RegFile[21][23]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux67~18_combout\)))) # (\R.curInst\(17) & ((!\Mux67~18_combout\ & ((\RegFile[22][23]~q\))) # (\Mux67~18_combout\ & (\RegFile[23][23]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][23]~q\,
	datab => \ALT_INV_RegFile[23][23]~q\,
	datac => \ALT_INV_RegFile[22][23]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux67~18_combout\,
	datag => \ALT_INV_RegFile[20][23]~q\,
	combout => \Mux67~5_combout\);

-- Location: LABCELL_X63_Y3_N36
\Decoder0~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~10_combout\ = ( !\R.curInst\(7) & ( \R.curInst\(9) & ( (\R.regWriteEn~q\ & (\R.curInst\(10) & (!\R.curInst\(11) & \R.curInst\(8)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000100000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.regWriteEn~q\,
	datab => \ALT_INV_R.curInst\(10),
	datac => \ALT_INV_R.curInst\(11),
	datad => \ALT_INV_R.curInst\(8),
	datae => \ALT_INV_R.curInst\(7),
	dataf => \ALT_INV_R.curInst\(9),
	combout => \Decoder0~10_combout\);

-- Location: FF_X62_Y2_N41
\RegFile[14][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(23),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][23]~q\);

-- Location: LABCELL_X64_Y5_N24
\Decoder0~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~7_combout\ = ( !\R.curInst\(8) & ( \R.curInst\(7) & ( (\R.curInst\(10) & (\R.regWriteEn~q\ & (!\R.curInst\(11) & \R.curInst\(9)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000100000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(10),
	datab => \ALT_INV_R.regWriteEn~q\,
	datac => \ALT_INV_R.curInst\(11),
	datad => \ALT_INV_R.curInst\(9),
	datae => \ALT_INV_R.curInst\(8),
	dataf => \ALT_INV_R.curInst\(7),
	combout => \Decoder0~7_combout\);

-- Location: FF_X62_Y2_N32
\RegFile[13][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(23),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][23]~q\);

-- Location: LABCELL_X63_Y3_N39
\Decoder0~20\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~20_combout\ = ( !\R.curInst\(9) & ( \R.curInst\(7) & ( (\R.regWriteEn~q\ & (\R.curInst\(10) & (\R.curInst\(8) & !\R.curInst\(11)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000001000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.regWriteEn~q\,
	datab => \ALT_INV_R.curInst\(10),
	datac => \ALT_INV_R.curInst\(8),
	datad => \ALT_INV_R.curInst\(11),
	datae => \ALT_INV_R.curInst\(9),
	dataf => \ALT_INV_R.curInst\(7),
	combout => \Decoder0~20_combout\);

-- Location: FF_X68_Y2_N44
\RegFile[11][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(23),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][23]~q\);

-- Location: LABCELL_X67_Y5_N15
\Decoder0~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~22_combout\ = ( \R.regWriteEn~q\ & ( !\R.curInst\(7) & ( (!\R.curInst\(11) & (\R.curInst\(10) & (\R.curInst\(8) & !\R.curInst\(9)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000100000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(11),
	datab => \ALT_INV_R.curInst\(10),
	datac => \ALT_INV_R.curInst\(8),
	datad => \ALT_INV_R.curInst\(9),
	datae => \ALT_INV_R.regWriteEn~q\,
	dataf => \ALT_INV_R.curInst\(7),
	combout => \Decoder0~22_combout\);

-- Location: FF_X59_Y3_N8
\RegFile[10][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(23),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][23]~q\);

-- Location: LABCELL_X68_Y5_N24
\Decoder0~19\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~19_combout\ = ( \R.curInst\(10) & ( !\R.curInst\(11) & ( (!\R.curInst\(9) & (!\R.curInst\(8) & (\R.curInst\(7) & \R.regWriteEn~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000100000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(9),
	datab => \ALT_INV_R.curInst\(8),
	datac => \ALT_INV_R.curInst\(7),
	datad => \ALT_INV_R.regWriteEn~q\,
	datae => \ALT_INV_R.curInst\(10),
	dataf => \ALT_INV_R.curInst\(11),
	combout => \Decoder0~19_combout\);

-- Location: FF_X68_Y2_N32
\RegFile[9][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(23),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][23]~q\);

-- Location: LABCELL_X66_Y5_N54
\RegFile[8][23]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[8][23]~feeder_combout\ = ( \R.regWriteData\(23) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(23),
	combout => \RegFile[8][23]~feeder_combout\);

-- Location: LABCELL_X68_Y5_N39
\Decoder0~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~21_combout\ = ( \R.curInst\(10) & ( !\R.curInst\(9) & ( (!\R.curInst\(11) & (!\R.curInst\(8) & (\R.regWriteEn~q\ & !\R.curInst\(7)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000010000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(11),
	datab => \ALT_INV_R.curInst\(8),
	datac => \ALT_INV_R.regWriteEn~q\,
	datad => \ALT_INV_R.curInst\(7),
	datae => \ALT_INV_R.curInst\(10),
	dataf => \ALT_INV_R.curInst\(9),
	combout => \Decoder0~21_combout\);

-- Location: FF_X66_Y5_N56
\RegFile[8][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[8][23]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][23]~q\);

-- Location: LABCELL_X68_Y2_N42
\Mux67~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux67~14_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & (\RegFile[8][23]~q\)) # (\R.curInst\(15) & ((\RegFile[9][23]~q\))))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & ((\RegFile[10][23]~q\))) # (\R.curInst\(15) & (\RegFile[11][23]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110000110011111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[11][23]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[10][23]~q\,
	datad => \ALT_INV_RegFile[9][23]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][23]~q\,
	combout => \Mux67~14_combout\);

-- Location: LABCELL_X63_Y3_N45
\Decoder0~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~9_combout\ = ( !\R.curInst\(8) & ( !\R.curInst\(11) & ( (\R.regWriteEn~q\ & (\R.curInst\(10) & (!\R.curInst\(7) & \R.curInst\(9)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000010000000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.regWriteEn~q\,
	datab => \ALT_INV_R.curInst\(10),
	datac => \ALT_INV_R.curInst\(7),
	datad => \ALT_INV_R.curInst\(9),
	datae => \ALT_INV_R.curInst\(8),
	dataf => \ALT_INV_R.curInst\(11),
	combout => \Decoder0~9_combout\);

-- Location: FF_X62_Y2_N43
\RegFile[12][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(23),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][23]~q\);

-- Location: LABCELL_X68_Y2_N54
\Mux67~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux67~1_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux67~14_combout\)))) # (\R.curInst\(17) & ((!\Mux67~14_combout\ & (\RegFile[12][23]~q\)) # (\Mux67~14_combout\ & ((\RegFile[13][23]~q\)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) 
-- & ((((\Mux67~14_combout\))))) # (\R.curInst\(17) & (((!\Mux67~14_combout\ & ((\RegFile[14][23]~q\))) # (\Mux67~14_combout\ & (\RegFile[15][23]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111001100111111111101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][23]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[14][23]~q\,
	datad => \ALT_INV_RegFile[13][23]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux67~14_combout\,
	datag => \ALT_INV_RegFile[12][23]~q\,
	combout => \Mux67~1_combout\);

-- Location: LABCELL_X67_Y5_N39
\Decoder0~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~6_combout\ = ( \R.regWriteEn~q\ & ( \R.curInst\(7) & ( (!\R.curInst\(11) & (\R.curInst\(8) & (!\R.curInst\(10) & !\R.curInst\(9)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000010000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(11),
	datab => \ALT_INV_R.curInst\(8),
	datac => \ALT_INV_R.curInst\(10),
	datad => \ALT_INV_R.curInst\(9),
	datae => \ALT_INV_R.regWriteEn~q\,
	dataf => \ALT_INV_R.curInst\(7),
	combout => \Decoder0~6_combout\);

-- Location: FF_X73_Y3_N14
\RegFile[3][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(23),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][23]~q\);

-- Location: LABCELL_X66_Y5_N3
\Decoder0~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~4_combout\ = ( !\R.curInst\(11) & ( \R.curInst\(8) & ( (!\R.curInst\(7) & (!\R.curInst\(9) & (\R.regWriteEn~q\ & !\R.curInst\(10)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000001000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(7),
	datab => \ALT_INV_R.curInst\(9),
	datac => \ALT_INV_R.regWriteEn~q\,
	datad => \ALT_INV_R.curInst\(10),
	datae => \ALT_INV_R.curInst\(11),
	dataf => \ALT_INV_R.curInst\(8),
	combout => \Decoder0~4_combout\);

-- Location: FF_X62_Y1_N8
\RegFile[2][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(23),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][23]~q\);

-- Location: LABCELL_X67_Y5_N9
\Decoder0~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~2_combout\ = ( \R.regWriteEn~q\ & ( !\R.curInst\(11) & ( (!\R.curInst\(7) & (!\R.curInst\(10) & (\R.curInst\(8) & \R.curInst\(9)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000100000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(7),
	datab => \ALT_INV_R.curInst\(10),
	datac => \ALT_INV_R.curInst\(8),
	datad => \ALT_INV_R.curInst\(9),
	datae => \ALT_INV_R.regWriteEn~q\,
	dataf => \ALT_INV_R.curInst\(11),
	combout => \Decoder0~2_combout\);

-- Location: FF_X73_Y3_N26
\RegFile[6][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(23),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][23]~q\);

-- Location: LABCELL_X68_Y5_N36
\Decoder0~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~0_combout\ = ( \R.curInst\(9) & ( !\R.curInst\(10) & ( (!\R.curInst\(11) & (!\R.curInst\(8) & (!\R.curInst\(7) & \R.regWriteEn~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000001000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(11),
	datab => \ALT_INV_R.curInst\(8),
	datac => \ALT_INV_R.curInst\(7),
	datad => \ALT_INV_R.regWriteEn~q\,
	datae => \ALT_INV_R.curInst\(9),
	dataf => \ALT_INV_R.curInst\(10),
	combout => \Decoder0~0_combout\);

-- Location: FF_X62_Y1_N55
\RegFile[4][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(23),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][23]~q\);

-- Location: LABCELL_X66_Y5_N30
\RegFile[5][23]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[5][23]~feeder_combout\ = ( \R.regWriteData\(23) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(23),
	combout => \RegFile[5][23]~feeder_combout\);

-- Location: LABCELL_X61_Y6_N39
\Decoder0~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~1_combout\ = ( \R.curInst\(7) & ( !\R.curInst\(8) & ( (\R.regWriteEn~q\ & (!\R.curInst\(11) & (\R.curInst\(9) & !\R.curInst\(10)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000001000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.regWriteEn~q\,
	datab => \ALT_INV_R.curInst\(11),
	datac => \ALT_INV_R.curInst\(9),
	datad => \ALT_INV_R.curInst\(10),
	datae => \ALT_INV_R.curInst\(7),
	dataf => \ALT_INV_R.curInst\(8),
	combout => \Decoder0~1_combout\);

-- Location: FF_X66_Y5_N31
\RegFile[5][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[5][23]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][23]~q\);

-- Location: LABCELL_X67_Y5_N33
\Decoder0~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~3_combout\ = ( \R.regWriteEn~q\ & ( \R.curInst\(9) & ( (!\R.curInst\(11) & (\R.curInst\(8) & (!\R.curInst\(10) & \R.curInst\(7)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000000000000100000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(11),
	datab => \ALT_INV_R.curInst\(8),
	datac => \ALT_INV_R.curInst\(10),
	datad => \ALT_INV_R.curInst\(7),
	datae => \ALT_INV_R.regWriteEn~q\,
	dataf => \ALT_INV_R.curInst\(9),
	combout => \Decoder0~3_combout\);

-- Location: FF_X73_Y3_N19
\RegFile[7][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(23),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][23]~q\);

-- Location: LABCELL_X73_Y3_N18
\Mux67~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux67~0_combout\ = ( \RegFile[7][23]~q\ & ( \R.curInst\(15) & ( (\R.curInst\(16)) # (\RegFile[5][23]~q\) ) ) ) # ( !\RegFile[7][23]~q\ & ( \R.curInst\(15) & ( (\RegFile[5][23]~q\ & !\R.curInst\(16)) ) ) ) # ( \RegFile[7][23]~q\ & ( !\R.curInst\(15) & ( 
-- (!\R.curInst\(16) & ((\RegFile[4][23]~q\))) # (\R.curInst\(16) & (\RegFile[6][23]~q\)) ) ) ) # ( !\RegFile[7][23]~q\ & ( !\R.curInst\(15) & ( (!\R.curInst\(16) & ((\RegFile[4][23]~q\))) # (\R.curInst\(16) & (\RegFile[6][23]~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001101010101001100110101010100001111000000000000111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[6][23]~q\,
	datab => \ALT_INV_RegFile[4][23]~q\,
	datac => \ALT_INV_RegFile[5][23]~q\,
	datad => \ALT_INV_R.curInst\(16),
	datae => \ALT_INV_RegFile[7][23]~q\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux67~0_combout\);

-- Location: LABCELL_X71_Y3_N6
\RegFile[1][23]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[1][23]~feeder_combout\ = ( \R.regWriteData\(23) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(23),
	combout => \RegFile[1][23]~feeder_combout\);

-- Location: LABCELL_X66_Y5_N12
\Decoder0~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~5_combout\ = ( !\R.curInst\(10) & ( !\R.curInst\(9) & ( (!\R.curInst\(11) & (\R.regWriteEn~q\ & (\R.curInst\(7) & !\R.curInst\(8)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001000000000000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(11),
	datab => \ALT_INV_R.regWriteEn~q\,
	datac => \ALT_INV_R.curInst\(7),
	datad => \ALT_INV_R.curInst\(8),
	datae => \ALT_INV_R.curInst\(10),
	dataf => \ALT_INV_R.curInst\(9),
	combout => \Decoder0~5_combout\);

-- Location: FF_X71_Y3_N7
\RegFile[1][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[1][23]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][23]~q\);

-- Location: LABCELL_X73_Y3_N12
\Mux67~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux67~26_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((\RegFile[1][23]~q\ & (\R.curInst\(15)))))) # (\R.curInst\(17) & ((((\Mux67~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & ((!\R.curInst\(15) & (((\RegFile[2][23]~q\)))) # 
-- (\R.curInst\(15) & (\RegFile[3][23]~q\)))) # (\R.curInst\(17) & ((((\Mux67~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001010000010100010001001010101010111110101111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[3][23]~q\,
	datac => \ALT_INV_RegFile[2][23]~q\,
	datad => \ALT_INV_R.curInst\(15),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux67~0_combout\,
	datag => \ALT_INV_RegFile[1][23]~q\,
	combout => \Mux67~26_combout\);

-- Location: LABCELL_X68_Y5_N3
\Decoder0~16\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~16_combout\ = ( \R.curInst\(7) & ( \R.curInst\(8) & ( (\R.curInst\(10) & (\R.curInst\(9) & (\R.regWriteEn~q\ & \R.curInst\(11)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000000000000000001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(10),
	datab => \ALT_INV_R.curInst\(9),
	datac => \ALT_INV_R.regWriteEn~q\,
	datad => \ALT_INV_R.curInst\(11),
	datae => \ALT_INV_R.curInst\(7),
	dataf => \ALT_INV_R.curInst\(8),
	combout => \Decoder0~16_combout\);

-- Location: FF_X70_Y3_N56
\RegFile[31][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(23),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][23]~q\);

-- Location: LABCELL_X68_Y5_N54
\Decoder0~15\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~15_combout\ = ( \R.curInst\(7) & ( !\R.curInst\(8) & ( (\R.curInst\(10) & (\R.curInst\(9) & (\R.curInst\(11) & \R.regWriteEn~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(10),
	datab => \ALT_INV_R.curInst\(9),
	datac => \ALT_INV_R.curInst\(11),
	datad => \ALT_INV_R.regWriteEn~q\,
	datae => \ALT_INV_R.curInst\(7),
	dataf => \ALT_INV_R.curInst\(8),
	combout => \Decoder0~15_combout\);

-- Location: FF_X63_Y2_N56
\RegFile[29][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(23),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][23]~q\);

-- Location: LABCELL_X66_Y3_N57
\RegFile[30][23]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[30][23]~feeder_combout\ = ( \R.regWriteData\(23) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(23),
	combout => \RegFile[30][23]~feeder_combout\);

-- Location: LABCELL_X68_Y5_N57
\Decoder0~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~18_combout\ = ( \R.curInst\(8) & ( !\R.curInst\(7) & ( (\R.curInst\(10) & (\R.curInst\(9) & (\R.regWriteEn~q\ & \R.curInst\(11)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(10),
	datab => \ALT_INV_R.curInst\(9),
	datac => \ALT_INV_R.regWriteEn~q\,
	datad => \ALT_INV_R.curInst\(11),
	datae => \ALT_INV_R.curInst\(8),
	dataf => \ALT_INV_R.curInst\(7),
	combout => \Decoder0~18_combout\);

-- Location: FF_X66_Y3_N58
\RegFile[30][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[30][23]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][23]~q\);

-- Location: LABCELL_X66_Y5_N51
\Decoder0~28\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~28_combout\ = ( \R.curInst\(11) & ( \R.curInst\(8) & ( (\R.curInst\(7) & (!\R.curInst\(9) & (\R.regWriteEn~q\ & \R.curInst\(10)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000000000000000100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(7),
	datab => \ALT_INV_R.curInst\(9),
	datac => \ALT_INV_R.regWriteEn~q\,
	datad => \ALT_INV_R.curInst\(10),
	datae => \ALT_INV_R.curInst\(11),
	dataf => \ALT_INV_R.curInst\(8),
	combout => \Decoder0~28_combout\);

-- Location: FF_X63_Y2_N32
\RegFile[27][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(23),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][23]~q\);

-- Location: LABCELL_X68_Y5_N6
\Decoder0~30\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~30_combout\ = ( \R.curInst\(10) & ( \R.curInst\(8) & ( (\R.curInst\(11) & (\R.regWriteEn~q\ & (!\R.curInst\(7) & !\R.curInst\(9)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000001000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(11),
	datab => \ALT_INV_R.regWriteEn~q\,
	datac => \ALT_INV_R.curInst\(7),
	datad => \ALT_INV_R.curInst\(9),
	datae => \ALT_INV_R.curInst\(10),
	dataf => \ALT_INV_R.curInst\(8),
	combout => \Decoder0~30_combout\);

-- Location: FF_X60_Y2_N37
\RegFile[26][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(23),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][23]~q\);

-- Location: LABCELL_X63_Y3_N9
\Decoder0~27\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~27_combout\ = ( \R.curInst\(10) & ( !\R.curInst\(8) & ( (\R.regWriteEn~q\ & (!\R.curInst\(9) & (\R.curInst\(7) & \R.curInst\(11)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000010000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.regWriteEn~q\,
	datab => \ALT_INV_R.curInst\(9),
	datac => \ALT_INV_R.curInst\(7),
	datad => \ALT_INV_R.curInst\(11),
	datae => \ALT_INV_R.curInst\(10),
	dataf => \ALT_INV_R.curInst\(8),
	combout => \Decoder0~27_combout\);

-- Location: FF_X63_Y2_N14
\RegFile[25][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(23),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][23]~q\);

-- Location: MLABCELL_X59_Y2_N6
\RegFile[24][23]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[24][23]~feeder_combout\ = ( \R.regWriteData\(23) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(23),
	combout => \RegFile[24][23]~feeder_combout\);

-- Location: LABCELL_X63_Y3_N33
\Decoder0~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~29_combout\ = ( \R.curInst\(10) & ( !\R.curInst\(8) & ( (\R.regWriteEn~q\ & (!\R.curInst\(7) & (\R.curInst\(11) & !\R.curInst\(9)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000001000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.regWriteEn~q\,
	datab => \ALT_INV_R.curInst\(7),
	datac => \ALT_INV_R.curInst\(11),
	datad => \ALT_INV_R.curInst\(9),
	datae => \ALT_INV_R.curInst\(10),
	dataf => \ALT_INV_R.curInst\(8),
	combout => \Decoder0~29_combout\);

-- Location: FF_X59_Y2_N7
\RegFile[24][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[24][23]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][23]~q\);

-- Location: LABCELL_X63_Y2_N30
\Mux67~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux67~22_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & (\RegFile[24][23]~q\)) # (\R.curInst\(15) & ((\RegFile[25][23]~q\)))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & ((\RegFile[26][23]~q\))) # (\R.curInst\(15) & (\RegFile[27][23]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001010101111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[27][23]~q\,
	datac => \ALT_INV_RegFile[26][23]~q\,
	datad => \ALT_INV_RegFile[25][23]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][23]~q\,
	combout => \Mux67~22_combout\);

-- Location: LABCELL_X73_Y2_N3
\RegFile[28][23]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[28][23]~feeder_combout\ = ( \R.regWriteData\(23) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(23),
	combout => \RegFile[28][23]~feeder_combout\);

-- Location: LABCELL_X67_Y6_N3
\Decoder0~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~17_combout\ = ( \R.curInst\(10) & ( !\R.curInst\(8) & ( (!\R.curInst\(7) & (\R.regWriteEn~q\ & (\R.curInst\(9) & \R.curInst\(11)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000001000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(7),
	datab => \ALT_INV_R.regWriteEn~q\,
	datac => \ALT_INV_R.curInst\(9),
	datad => \ALT_INV_R.curInst\(11),
	datae => \ALT_INV_R.curInst\(10),
	dataf => \ALT_INV_R.curInst\(8),
	combout => \Decoder0~17_combout\);

-- Location: FF_X73_Y2_N4
\RegFile[28][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[28][23]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][23]~q\);

-- Location: LABCELL_X70_Y3_N54
\Mux67~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux67~9_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux67~22_combout\)))) # (\R.curInst\(17) & ((!\Mux67~22_combout\ & ((\RegFile[28][23]~q\))) # (\Mux67~22_combout\ & (\RegFile[29][23]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux67~22_combout\)))) # (\R.curInst\(17) & ((!\Mux67~22_combout\ & ((\RegFile[30][23]~q\))) # (\Mux67~22_combout\ & (\RegFile[31][23]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][23]~q\,
	datab => \ALT_INV_RegFile[29][23]~q\,
	datac => \ALT_INV_RegFile[30][23]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux67~22_combout\,
	datag => \ALT_INV_RegFile[28][23]~q\,
	combout => \Mux67~9_combout\);

-- Location: LABCELL_X71_Y3_N36
\Mux67~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux67~13_combout\ = ( \Mux67~26_combout\ & ( \Mux67~9_combout\ & ( (!\R.curInst\(18) & ((!\R.curInst\(19)) # ((\Mux67~5_combout\)))) # (\R.curInst\(18) & (((\Mux67~1_combout\)) # (\R.curInst\(19)))) ) ) ) # ( !\Mux67~26_combout\ & ( \Mux67~9_combout\ & ( 
-- (!\R.curInst\(18) & (\R.curInst\(19) & (\Mux67~5_combout\))) # (\R.curInst\(18) & (((\Mux67~1_combout\)) # (\R.curInst\(19)))) ) ) ) # ( \Mux67~26_combout\ & ( !\Mux67~9_combout\ & ( (!\R.curInst\(18) & ((!\R.curInst\(19)) # ((\Mux67~5_combout\)))) # 
-- (\R.curInst\(18) & (!\R.curInst\(19) & ((\Mux67~1_combout\)))) ) ) ) # ( !\Mux67~26_combout\ & ( !\Mux67~9_combout\ & ( (!\R.curInst\(18) & (\R.curInst\(19) & (\Mux67~5_combout\))) # (\R.curInst\(18) & (!\R.curInst\(19) & ((\Mux67~1_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001001000110100010101100111000010011010101111001101111011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(18),
	datab => \ALT_INV_R.curInst\(19),
	datac => \ALT_INV_Mux67~5_combout\,
	datad => \ALT_INV_Mux67~1_combout\,
	datae => \ALT_INV_Mux67~26_combout\,
	dataf => \ALT_INV_Mux67~9_combout\,
	combout => \Mux67~13_combout\);

-- Location: LABCELL_X74_Y3_N18
\Mux231~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux231~0_combout\ = ( \Mux67~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC\(23)))) ) ) # ( !\Mux67~13_combout\ & ( (\vAluSrc1~2_combout\ & (\R.curPC\(23) & !\vAluSrc1~1_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000000000000110000000011001111000000001100111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_vAluSrc1~2_combout\,
	datac => \ALT_INV_R.curPC\(23),
	datad => \ALT_INV_vAluSrc1~1_combout\,
	dataf => \ALT_INV_Mux67~13_combout\,
	combout => \Mux231~0_combout\);

-- Location: FF_X74_Y3_N16
\R.aluData1[23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux231~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData1\(23));

-- Location: LABCELL_X74_Y4_N45
\Mux132~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux132~0_combout\ = ( \Mux123~1_combout\ ) # ( !\Mux123~1_combout\ & ( (\vAluSrc1~0_combout\ & (((\R.curInst\(2) & \R.curInst\(22))) # (\Mux124~0_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000111000001010000011111111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux124~0_combout\,
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_vAluSrc1~0_combout\,
	datad => \ALT_INV_R.curInst\(22),
	dataf => \ALT_INV_Mux123~1_combout\,
	combout => \Mux132~0_combout\);

-- Location: LABCELL_X77_Y5_N6
\Equal4~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Equal4~0_combout\ = ( \R.curInst\(5) & ( (\R.curInst\(2) & (!\R.curInst\(4) & \R.curInst\(6))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000010001000000000001000100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(2),
	datab => \ALT_INV_R.curInst\(4),
	datad => \ALT_INV_R.curInst\(6),
	dataf => \ALT_INV_R.curInst\(5),
	combout => \Equal4~0_combout\);

-- Location: MLABCELL_X78_Y4_N27
\Equal4~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Equal4~2_combout\ = ( \Equal4~0_combout\ & ( (!\R.curInst\(3) & \Equal4~1_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000111100000000000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.curInst\(3),
	datad => \ALT_INV_Equal4~1_combout\,
	dataf => \ALT_INV_Equal4~0_combout\,
	combout => \Equal4~2_combout\);

-- Location: FF_X64_Y1_N44
\RegFile[21][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(22),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][22]~q\);

-- Location: FF_X70_Y3_N26
\RegFile[23][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(22),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][22]~q\);

-- Location: FF_X59_Y4_N43
\RegFile[22][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(22),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][22]~q\);

-- Location: FF_X64_Y1_N8
\RegFile[17][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(22),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][22]~q\);

-- Location: FF_X70_Y3_N44
\RegFile[19][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(22),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][22]~q\);

-- Location: MLABCELL_X59_Y3_N36
\RegFile[18][22]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[18][22]~feeder_combout\ = ( \R.regWriteData\(22) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(22),
	combout => \RegFile[18][22]~feeder_combout\);

-- Location: FF_X59_Y3_N37
\RegFile[18][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][22]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][22]~q\);

-- Location: LABCELL_X64_Y1_N18
\RegFile[16][22]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[16][22]~feeder_combout\ = ( \R.regWriteData\(22) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(22),
	combout => \RegFile[16][22]~feeder_combout\);

-- Location: FF_X64_Y1_N19
\RegFile[16][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[16][22]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][22]~q\);

-- Location: LABCELL_X70_Y3_N42
\Mux68~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux68~18_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[16][22]~q\))) # (\R.curInst\(15) & (\RegFile[17][22]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[18][22]~q\))) # (\R.curInst\(15) & (\RegFile[19][22]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[17][22]~q\,
	datab => \ALT_INV_RegFile[19][22]~q\,
	datac => \ALT_INV_RegFile[18][22]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][22]~q\,
	combout => \Mux68~18_combout\);

-- Location: FF_X59_Y4_N58
\RegFile[20][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(22),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][22]~q\);

-- Location: LABCELL_X70_Y3_N24
\Mux68~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux68~5_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux68~18_combout\)))) # (\R.curInst\(17) & ((!\Mux68~18_combout\ & ((\RegFile[20][22]~q\))) # (\Mux68~18_combout\ & (\RegFile[21][22]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux68~18_combout\)))) # (\R.curInst\(17) & ((!\Mux68~18_combout\ & ((\RegFile[22][22]~q\))) # (\Mux68~18_combout\ & (\RegFile[23][22]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][22]~q\,
	datab => \ALT_INV_RegFile[23][22]~q\,
	datac => \ALT_INV_RegFile[22][22]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux68~18_combout\,
	datag => \ALT_INV_RegFile[20][22]~q\,
	combout => \Mux68~5_combout\);

-- Location: FF_X73_Y2_N7
\RegFile[30][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(22),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][22]~q\);

-- Location: FF_X63_Y2_N26
\RegFile[29][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(22),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][22]~q\);

-- Location: FF_X63_Y2_N38
\RegFile[27][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(22),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][22]~q\);

-- Location: FF_X63_Y2_N20
\RegFile[25][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(22),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][22]~q\);

-- Location: LABCELL_X60_Y2_N30
\RegFile[26][22]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[26][22]~feeder_combout\ = ( \R.regWriteData\(22) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(22),
	combout => \RegFile[26][22]~feeder_combout\);

-- Location: FF_X60_Y2_N31
\RegFile[26][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[26][22]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][22]~q\);

-- Location: MLABCELL_X59_Y2_N12
\RegFile[24][22]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[24][22]~feeder_combout\ = ( \R.regWriteData\(22) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(22),
	combout => \RegFile[24][22]~feeder_combout\);

-- Location: FF_X59_Y2_N13
\RegFile[24][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[24][22]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][22]~q\);

-- Location: LABCELL_X63_Y2_N36
\Mux68~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux68~22_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[24][22]~q\))) # (\R.curInst\(15) & (\RegFile[25][22]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[26][22]~q\))) # (\R.curInst\(15) & (\RegFile[27][22]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[27][22]~q\,
	datab => \ALT_INV_RegFile[25][22]~q\,
	datac => \ALT_INV_RegFile[26][22]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][22]~q\,
	combout => \Mux68~22_combout\);

-- Location: FF_X73_Y2_N31
\RegFile[28][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(22),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][22]~q\);

-- Location: LABCELL_X70_Y3_N30
\Mux68~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux68~9_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux68~22_combout\))))) # (\R.curInst\(17) & (((!\Mux68~22_combout\ & (\RegFile[28][22]~q\)) # (\Mux68~22_combout\ & ((\RegFile[29][22]~q\)))))) ) ) # ( \R.curInst\(16) & ( 
-- (!\R.curInst\(17) & ((((\Mux68~22_combout\))))) # (\R.curInst\(17) & (((!\Mux68~22_combout\ & ((\RegFile[30][22]~q\))) # (\Mux68~22_combout\ & (\RegFile[31][22]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110101010111111111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[31][22]~q\,
	datac => \ALT_INV_RegFile[30][22]~q\,
	datad => \ALT_INV_RegFile[29][22]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux68~22_combout\,
	datag => \ALT_INV_RegFile[28][22]~q\,
	combout => \Mux68~9_combout\);

-- Location: FF_X68_Y3_N56
\RegFile[3][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(22),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][22]~q\);

-- Location: FF_X62_Y1_N50
\RegFile[2][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(22),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][22]~q\);

-- Location: LABCELL_X62_Y1_N27
\RegFile[4][22]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[4][22]~feeder_combout\ = ( \R.regWriteData\(22) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(22),
	combout => \RegFile[4][22]~feeder_combout\);

-- Location: FF_X62_Y1_N28
\RegFile[4][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[4][22]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][22]~q\);

-- Location: FF_X68_Y3_N37
\RegFile[5][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(22),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][22]~q\);

-- Location: FF_X59_Y5_N28
\RegFile[6][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(22),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][22]~q\);

-- Location: FF_X68_Y3_N19
\RegFile[7][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(22),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][22]~q\);

-- Location: LABCELL_X68_Y3_N18
\Mux68~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux68~0_combout\ = ( \RegFile[7][22]~q\ & ( \R.curInst\(15) & ( (\R.curInst\(16)) # (\RegFile[5][22]~q\) ) ) ) # ( !\RegFile[7][22]~q\ & ( \R.curInst\(15) & ( (\RegFile[5][22]~q\ & !\R.curInst\(16)) ) ) ) # ( \RegFile[7][22]~q\ & ( !\R.curInst\(15) & ( 
-- (!\R.curInst\(16) & (\RegFile[4][22]~q\)) # (\R.curInst\(16) & ((\RegFile[6][22]~q\))) ) ) ) # ( !\RegFile[7][22]~q\ & ( !\R.curInst\(15) & ( (!\R.curInst\(16) & (\RegFile[4][22]~q\)) # (\R.curInst\(16) & ((\RegFile[6][22]~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010100001111010101010000111100110011000000000011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[4][22]~q\,
	datab => \ALT_INV_RegFile[5][22]~q\,
	datac => \ALT_INV_RegFile[6][22]~q\,
	datad => \ALT_INV_R.curInst\(16),
	datae => \ALT_INV_RegFile[7][22]~q\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux68~0_combout\);

-- Location: MLABCELL_X72_Y3_N39
\RegFile[1][22]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[1][22]~feeder_combout\ = \R.regWriteData\(22)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.regWriteData\(22),
	combout => \RegFile[1][22]~feeder_combout\);

-- Location: FF_X72_Y3_N41
\RegFile[1][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[1][22]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][22]~q\);

-- Location: LABCELL_X68_Y3_N54
\Mux68~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux68~26_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (\RegFile[1][22]~q\ & (\R.curInst\(15)))) # (\R.curInst\(17) & (((\Mux68~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & ((!\R.curInst\(15) & (((\RegFile[2][22]~q\)))) # 
-- (\R.curInst\(15) & (\RegFile[3][22]~q\)))) # (\R.curInst\(17) & ((((\Mux68~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001100000011000100010000110011001111110011111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][22]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[2][22]~q\,
	datad => \ALT_INV_R.curInst\(15),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux68~0_combout\,
	datag => \ALT_INV_RegFile[1][22]~q\,
	combout => \Mux68~26_combout\);

-- Location: FF_X62_Y2_N2
\RegFile[13][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(22),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][22]~q\);

-- Location: LABCELL_X62_Y2_N36
\RegFile[14][22]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[14][22]~feeder_combout\ = \R.regWriteData\(22)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110011001100110011001100110011001100110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.regWriteData\(22),
	combout => \RegFile[14][22]~feeder_combout\);

-- Location: FF_X62_Y2_N38
\RegFile[14][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[14][22]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][22]~q\);

-- Location: LABCELL_X63_Y3_N3
\Decoder0~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \Decoder0~8_combout\ = ( \R.curInst\(8) & ( \R.curInst\(7) & ( (\R.regWriteEn~q\ & (\R.curInst\(9) & (\R.curInst\(10) & !\R.curInst\(11)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000000000100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.regWriteEn~q\,
	datab => \ALT_INV_R.curInst\(9),
	datac => \ALT_INV_R.curInst\(10),
	datad => \ALT_INV_R.curInst\(11),
	datae => \ALT_INV_R.curInst\(8),
	dataf => \ALT_INV_R.curInst\(7),
	combout => \Decoder0~8_combout\);

-- Location: FF_X68_Y2_N2
\RegFile[15][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(22),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][22]~q\);

-- Location: FF_X68_Y2_N26
\RegFile[11][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(22),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][22]~q\);

-- Location: MLABCELL_X59_Y3_N33
\RegFile[10][22]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[10][22]~feeder_combout\ = ( \R.regWriteData\(22) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(22),
	combout => \RegFile[10][22]~feeder_combout\);

-- Location: FF_X59_Y3_N34
\RegFile[10][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[10][22]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][22]~q\);

-- Location: FF_X68_Y2_N14
\RegFile[9][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(22),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][22]~q\);

-- Location: FF_X68_Y5_N1
\RegFile[8][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(22),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][22]~q\);

-- Location: LABCELL_X68_Y2_N24
\Mux68~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux68~14_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & (\RegFile[8][22]~q\)) # (\R.curInst\(15) & ((\RegFile[9][22]~q\)))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & ((\RegFile[10][22]~q\))) # (\R.curInst\(15) & (\RegFile[11][22]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001010101111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[11][22]~q\,
	datac => \ALT_INV_RegFile[10][22]~q\,
	datad => \ALT_INV_RegFile[9][22]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][22]~q\,
	combout => \Mux68~14_combout\);

-- Location: LABCELL_X62_Y2_N9
\RegFile[12][22]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[12][22]~feeder_combout\ = \R.regWriteData\(22)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.regWriteData\(22),
	combout => \RegFile[12][22]~feeder_combout\);

-- Location: FF_X62_Y2_N11
\RegFile[12][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[12][22]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][22]~q\);

-- Location: LABCELL_X68_Y2_N0
\Mux68~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux68~1_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux68~14_combout\))))) # (\R.curInst\(17) & (((!\Mux68~14_combout\ & ((\RegFile[12][22]~q\))) # (\Mux68~14_combout\ & (\RegFile[13][22]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- (!\R.curInst\(17) & ((((\Mux68~14_combout\))))) # (\R.curInst\(17) & (((!\Mux68~14_combout\ & (\RegFile[14][22]~q\)) # (\Mux68~14_combout\ & ((\RegFile[15][22]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110111011101110111010101011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[13][22]~q\,
	datac => \ALT_INV_RegFile[14][22]~q\,
	datad => \ALT_INV_RegFile[15][22]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux68~14_combout\,
	datag => \ALT_INV_RegFile[12][22]~q\,
	combout => \Mux68~1_combout\);

-- Location: LABCELL_X70_Y3_N36
\Mux68~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux68~13_combout\ = ( \Mux68~26_combout\ & ( \Mux68~1_combout\ & ( (!\R.curInst\(19)) # ((!\R.curInst\(18) & (\Mux68~5_combout\)) # (\R.curInst\(18) & ((\Mux68~9_combout\)))) ) ) ) # ( !\Mux68~26_combout\ & ( \Mux68~1_combout\ & ( (!\R.curInst\(18) & 
-- (\R.curInst\(19) & (\Mux68~5_combout\))) # (\R.curInst\(18) & ((!\R.curInst\(19)) # ((\Mux68~9_combout\)))) ) ) ) # ( \Mux68~26_combout\ & ( !\Mux68~1_combout\ & ( (!\R.curInst\(18) & ((!\R.curInst\(19)) # ((\Mux68~5_combout\)))) # (\R.curInst\(18) & 
-- (\R.curInst\(19) & ((\Mux68~9_combout\)))) ) ) ) # ( !\Mux68~26_combout\ & ( !\Mux68~1_combout\ & ( (\R.curInst\(19) & ((!\R.curInst\(18) & (\Mux68~5_combout\)) # (\R.curInst\(18) & ((\Mux68~9_combout\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001000010011100010101001101101000110010101111100111011011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(18),
	datab => \ALT_INV_R.curInst\(19),
	datac => \ALT_INV_Mux68~5_combout\,
	datad => \ALT_INV_Mux68~9_combout\,
	datae => \ALT_INV_Mux68~26_combout\,
	dataf => \ALT_INV_Mux68~1_combout\,
	combout => \Mux68~13_combout\);

-- Location: LABCELL_X74_Y3_N48
\Mux232~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux232~0_combout\ = ( \Mux68~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC\(22)))) ) ) # ( !\Mux68~13_combout\ & ( (\vAluSrc1~2_combout\ & (\R.curPC\(22) & !\vAluSrc1~1_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000000000000110000000011001111000000001100111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_vAluSrc1~2_combout\,
	datac => \ALT_INV_R.curPC\(22),
	datad => \ALT_INV_vAluSrc1~1_combout\,
	dataf => \ALT_INV_Mux68~13_combout\,
	combout => \Mux232~0_combout\);

-- Location: FF_X74_Y3_N47
\R.aluData1[22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux232~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData1\(22));

-- Location: FF_X71_Y7_N5
\R.aluOp.ALUOpSLL\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.aluOp.ALUOpSLL_OTERM359\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluOp.ALUOpSLL~q\);

-- Location: LABCELL_X77_Y3_N9
\Mux26~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux26~0_combout\ = ( \R.curInst\(5) & ( (!\R.curInst\(2)) # (\R.curInst\(6)) ) ) # ( !\R.curInst\(5) & ( (!\R.curInst\(2) & !\R.curInst\(6)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010101000000000101010100000000010101010111111111010101011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(2),
	datad => \ALT_INV_R.curInst\(6),
	dataf => \ALT_INV_R.curInst\(5),
	combout => \Mux26~0_combout\);

-- Location: LABCELL_X77_Y6_N27
\Mux162~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux162~0_combout\ = ( !\R.curInst\(13) & ( \R.curInst\(12) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111000000001111111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \ALT_INV_R.curInst\(12),
	dataf => \ALT_INV_R.curInst\(13),
	combout => \Mux162~0_combout\);

-- Location: LABCELL_X77_Y6_N33
\Mux24~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux24~0_combout\ = ( \Mux162~0_combout\ & ( (!\R.curInst\(6) & (!\R.curInst\(2) & (!\R.curInst\(14)))) # (\R.curInst\(6) & (((\R.aluOp.ALUOpSLL~q\)))) ) ) # ( !\Mux162~0_combout\ & ( (\R.curInst\(6) & \R.aluOp.ALUOpSLL~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010101000000000101010110000000110101011000000011010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(6),
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_R.curInst\(14),
	datad => \ALT_INV_R.aluOp.ALUOpSLL~q\,
	dataf => \ALT_INV_Mux162~0_combout\,
	combout => \Mux24~0_combout\);

-- Location: LABCELL_X77_Y6_N54
\Mux24~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux24~1_combout\ = ( \R.aluOp.ALUOpSLL~q\ & ( \Mux24~0_combout\ & ( ((!\R.curInst\(3) & (!\Mux26~0_combout\)) # (\R.curInst\(3) & ((!\Mux123~0_combout\)))) # (\R.curInst\(4)) ) ) ) # ( !\R.aluOp.ALUOpSLL~q\ & ( \Mux24~0_combout\ & ( (!\R.curInst\(3) & 
-- \R.curInst\(4)) ) ) ) # ( \R.aluOp.ALUOpSLL~q\ & ( !\Mux24~0_combout\ & ( (!\R.curInst\(3) & (!\Mux26~0_combout\ & (!\R.curInst\(4)))) # (\R.curInst\(3) & (((!\Mux123~0_combout\) # (\R.curInst\(4))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110101011000010100001010000010101101111110001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(3),
	datab => \ALT_INV_Mux26~0_combout\,
	datac => \ALT_INV_R.curInst\(4),
	datad => \ALT_INV_Mux123~0_combout\,
	datae => \ALT_INV_R.aluOp.ALUOpSLL~q\,
	dataf => \ALT_INV_Mux24~0_combout\,
	combout => \Mux24~1_combout\);

-- Location: LABCELL_X71_Y7_N33
\R.aluOp.ALUOpSLL_NEW358\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.aluOp.ALUOpSLL_OTERM359\ = ( \Mux24~1_combout\ & ( (\R.aluOp.ALUOpSLL~q\) # (\vAluSrc2~0_combout\) ) ) # ( !\Mux24~1_combout\ & ( (!\vAluSrc2~0_combout\ & \R.aluOp.ALUOpSLL~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011110000000000001111000000001111111111110000111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_vAluSrc2~0_combout\,
	datad => \ALT_INV_R.aluOp.ALUOpSLL~q\,
	dataf => \ALT_INV_Mux24~1_combout\,
	combout => \R.aluOp.ALUOpSLL_OTERM359\);

-- Location: LABCELL_X77_Y5_N21
\Mux150~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux150~0_combout\ = ( \R.curInst\(11) & ( \R.curInst\(24) & ( ((\Mux53~0_combout\ & ((\Mux18~0_combout\) # (\Mux154~0_combout\)))) # (\Equal4~0_combout\) ) ) ) # ( !\R.curInst\(11) & ( \R.curInst\(24) & ( ((\Mux53~0_combout\ & \Mux154~0_combout\)) # 
-- (\Equal4~0_combout\) ) ) ) # ( \R.curInst\(11) & ( !\R.curInst\(24) & ( (\Mux53~0_combout\ & \Mux18~0_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000001010000010100010001111111110001010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux53~0_combout\,
	datab => \ALT_INV_Mux154~0_combout\,
	datac => \ALT_INV_Mux18~0_combout\,
	datad => \ALT_INV_Equal4~0_combout\,
	datae => \ALT_INV_R.curInst\(11),
	dataf => \ALT_INV_R.curInst\(24),
	combout => \Mux150~0_combout\);

-- Location: FF_X77_Y6_N38
\R.aluOp.ALUOpSRL\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \R.aluOp.ALUOpSRL_OTERM361\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluOp.ALUOpSRL~q\);

-- Location: LABCELL_X77_Y6_N3
\Mux21~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux21~0_combout\ = ( !\R.curInst\(2) & ( (\R.curInst\(14) & !\R.curInst\(6)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100000000000011110000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.curInst\(14),
	datad => \ALT_INV_R.curInst\(6),
	dataf => \ALT_INV_R.curInst\(2),
	combout => \Mux21~0_combout\);

-- Location: LABCELL_X77_Y6_N12
\Mux25~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux25~0_combout\ = ( \Mux162~0_combout\ & ( (!\Mux21~0_combout\ & (\R.curInst\(6) & (\R.aluOp.ALUOpSRL~q\))) # (\Mux21~0_combout\ & ((!\R.curInst\(30)) # ((\R.curInst\(6) & \R.aluOp.ALUOpSRL~q\)))) ) ) # ( !\Mux162~0_combout\ & ( (\R.curInst\(6) & 
-- \R.aluOp.ALUOpSRL~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000110000001101010111000000110101011100000011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux21~0_combout\,
	datab => \ALT_INV_R.curInst\(6),
	datac => \ALT_INV_R.aluOp.ALUOpSRL~q\,
	datad => \ALT_INV_R.curInst\(30),
	dataf => \ALT_INV_Mux162~0_combout\,
	combout => \Mux25~0_combout\);

-- Location: LABCELL_X77_Y6_N42
\Mux25~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux25~1_combout\ = ( \R.aluOp.ALUOpSRL~q\ & ( \Mux25~0_combout\ & ( ((!\R.curInst\(3) & (!\Mux26~0_combout\)) # (\R.curInst\(3) & ((!\Mux123~0_combout\)))) # (\R.curInst\(4)) ) ) ) # ( !\R.aluOp.ALUOpSRL~q\ & ( \Mux25~0_combout\ & ( (\R.curInst\(4) & 
-- !\R.curInst\(3)) ) ) ) # ( \R.aluOp.ALUOpSRL~q\ & ( !\Mux25~0_combout\ & ( (!\R.curInst\(4) & ((!\R.curInst\(3) & (!\Mux26~0_combout\)) # (\R.curInst\(3) & ((!\Mux123~0_combout\))))) # (\R.curInst\(4) & (((\R.curInst\(3))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000100011111000010101010000010100001101111111010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(4),
	datab => \ALT_INV_Mux26~0_combout\,
	datac => \ALT_INV_R.curInst\(3),
	datad => \ALT_INV_Mux123~0_combout\,
	datae => \ALT_INV_R.aluOp.ALUOpSRL~q\,
	dataf => \ALT_INV_Mux25~0_combout\,
	combout => \Mux25~1_combout\);

-- Location: LABCELL_X77_Y6_N36
\R.aluOp.ALUOpSRL_NEW360\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.aluOp.ALUOpSRL_OTERM361\ = ( \vAluSrc2~0_combout\ & ( \Mux25~1_combout\ ) ) # ( !\vAluSrc2~0_combout\ & ( \R.aluOp.ALUOpSRL~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111000000001111111100110011001100110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Mux25~1_combout\,
	datad => \ALT_INV_R.aluOp.ALUOpSRL~q\,
	dataf => \ALT_INV_vAluSrc2~0_combout\,
	combout => \R.aluOp.ALUOpSRL_OTERM361\);

-- Location: MLABCELL_X72_Y5_N24
\Selector31~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector31~7_combout\ = (\R.aluOp.ALUOpSRL_OTERM361\ & \NxR.aluData2[4]~20_combout\)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000001111000000000000111100000000000011110000000000001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluOp.ALUOpSRL_OTERM361\,
	datad => \ALT_INV_NxR.aluData2[4]~20_combout\,
	combout => \Selector31~7_combout\);

-- Location: FF_X72_Y5_N25
\Selector31~7_NEW_REG382\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector31~7_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector31~7_OTERM383\);

-- Location: FF_X77_Y6_N41
\Selector31~0_NEW_REG348\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector31~0_NEW_REG348_OTERM569\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector31~0_OTERM349\);

-- Location: LABCELL_X77_Y6_N30
\R.aluOp.ALUOpSRA_NEW362\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.aluOp.ALUOpSRA_OTERM363\ = ( \vAluSrc2~0_combout\ & ( \Mux26~2_combout\ ) ) # ( !\vAluSrc2~0_combout\ & ( \R.aluOp.ALUOpSRA~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111000000001111111100001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Mux26~2_combout\,
	datad => \ALT_INV_R.aluOp.ALUOpSRA~q\,
	dataf => \ALT_INV_vAluSrc2~0_combout\,
	combout => \R.aluOp.ALUOpSRA_OTERM363\);

-- Location: FF_X77_Y6_N32
\R.aluOp.ALUOpSRA\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \R.aluOp.ALUOpSRA_OTERM363\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluOp.ALUOpSRA~q\);

-- Location: LABCELL_X77_Y6_N24
\Mux26~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux26~1_combout\ = ( \Mux162~0_combout\ & ( (!\R.curInst\(30) & (\R.curInst\(6) & ((\R.aluOp.ALUOpSRA~q\)))) # (\R.curInst\(30) & (((\R.curInst\(6) & \R.aluOp.ALUOpSRA~q\)) # (\Mux21~0_combout\))) ) ) # ( !\Mux162~0_combout\ & ( (\R.curInst\(6) & 
-- \R.aluOp.ALUOpSRA~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110011000000000011001100000101001101110000010100110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(30),
	datab => \ALT_INV_R.curInst\(6),
	datac => \ALT_INV_Mux21~0_combout\,
	datad => \ALT_INV_R.aluOp.ALUOpSRA~q\,
	dataf => \ALT_INV_Mux162~0_combout\,
	combout => \Mux26~1_combout\);

-- Location: LABCELL_X77_Y6_N51
\Mux26~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux26~2_combout\ = ( \R.aluOp.ALUOpSRA~q\ & ( \Mux26~1_combout\ & ( ((!\R.curInst\(3) & (!\Mux26~0_combout\)) # (\R.curInst\(3) & ((!\Mux123~0_combout\)))) # (\R.curInst\(4)) ) ) ) # ( !\R.aluOp.ALUOpSRA~q\ & ( \Mux26~1_combout\ & ( (\R.curInst\(4) & 
-- !\R.curInst\(3)) ) ) ) # ( \R.aluOp.ALUOpSRA~q\ & ( !\Mux26~1_combout\ & ( (!\R.curInst\(4) & ((!\R.curInst\(3) & (!\Mux26~0_combout\)) # (\R.curInst\(3) & ((!\Mux123~0_combout\))))) # (\R.curInst\(4) & (((\R.curInst\(3))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000100010001111010101010101000000001101110111110101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(4),
	datab => \ALT_INV_Mux26~0_combout\,
	datac => \ALT_INV_Mux123~0_combout\,
	datad => \ALT_INV_R.curInst\(3),
	datae => \ALT_INV_R.aluOp.ALUOpSRA~q\,
	dataf => \ALT_INV_Mux26~1_combout\,
	combout => \Mux26~2_combout\);

-- Location: LABCELL_X77_Y6_N39
\Selector31~0_NEW_REG348_NEW568\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector31~0_NEW_REG348_OTERM569\ = ( \Mux26~2_combout\ & ( (\Selector31~0_OTERM349\) # (\vAluSrc2~0_combout\) ) ) # ( !\Mux26~2_combout\ & ( (!\vAluSrc2~0_combout\ & ((\Selector31~0_OTERM349\))) # (\vAluSrc2~0_combout\ & (\Mux25~1_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000110111011000100011011101101010101111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluSrc2~0_combout\,
	datab => \ALT_INV_Mux25~1_combout\,
	datad => \ALT_INV_Selector31~0_OTERM349\,
	dataf => \ALT_INV_Mux26~2_combout\,
	combout => \Selector31~0_NEW_REG348_OTERM569\);

-- Location: LABCELL_X77_Y6_N18
\Selector31~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector31~5_combout\ = ( !\NxR.aluData2[4]~20_combout\ & ( \Selector31~0_NEW_REG348_OTERM569\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111000000001111111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \ALT_INV_Selector31~0_NEW_REG348_OTERM569\,
	dataf => \ALT_INV_NxR.aluData2[4]~20_combout\,
	combout => \Selector31~5_combout\);

-- Location: FF_X77_Y6_N19
\Selector31~5_NEW_REG598\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector31~5_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector31~5_OTERM599\);

-- Location: LABCELL_X77_Y5_N3
\Mux152~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux152~0_combout\ = ( \R.curInst\(22) & ( \R.curInst\(9) & ( ((\Mux53~0_combout\ & ((\Mux18~0_combout\) # (\Mux154~0_combout\)))) # (\Equal4~0_combout\) ) ) ) # ( !\R.curInst\(22) & ( \R.curInst\(9) & ( (\Mux53~0_combout\ & \Mux18~0_combout\) ) ) ) # ( 
-- \R.curInst\(22) & ( !\R.curInst\(9) & ( ((\Mux53~0_combout\ & \Mux154~0_combout\)) # (\Equal4~0_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000100011111111100000101000001010001010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux53~0_combout\,
	datab => \ALT_INV_Mux154~0_combout\,
	datac => \ALT_INV_Mux18~0_combout\,
	datad => \ALT_INV_Equal4~0_combout\,
	datae => \ALT_INV_R.curInst\(22),
	dataf => \ALT_INV_R.curInst\(9),
	combout => \Mux152~0_combout\);

-- Location: MLABCELL_X72_Y5_N51
\Selector31~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector31~6_combout\ = ( \R.aluOp.ALUOpSRA_OTERM363\ & ( \NxR.aluData2[4]~20_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000111111110000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \ALT_INV_NxR.aluData2[4]~20_combout\,
	dataf => \ALT_INV_R.aluOp.ALUOpSRA_OTERM363\,
	combout => \Selector31~6_combout\);

-- Location: FF_X72_Y5_N52
\Selector31~6_NEW_REG380\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector31~6_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector31~6_OTERM381\);

-- Location: FF_X71_Y7_N46
\R.aluData2[2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \NxR.aluData2[2]~19_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData2\(2));

-- Location: FF_X73_Y5_N16
\R.aluData1[28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux226~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData1\(28));

-- Location: LABCELL_X74_Y4_N0
\Mux127~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux127~0_combout\ = ( \Mux124~0_combout\ & ( (\Mux123~1_combout\) # (\vAluSrc1~0_combout\) ) ) # ( !\Mux124~0_combout\ & ( ((\vAluSrc1~0_combout\ & (\R.curInst\(2) & \R.curInst\(27)))) # (\Mux123~1_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000111111111000000011111111101010101111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluSrc1~0_combout\,
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_R.curInst\(27),
	datad => \ALT_INV_Mux123~1_combout\,
	dataf => \ALT_INV_Mux124~0_combout\,
	combout => \Mux127~0_combout\);

-- Location: LABCELL_X74_Y4_N15
\Mux123~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux123~3_combout\ = ( \R.curInst\(5) & ( ((\R.curInst\(31) & (\R.curInst\(2) & \vAluSrc1~0_combout\))) # (\Mux123~1_combout\) ) ) # ( !\R.curInst\(5) & ( ((\R.curInst\(31) & \vAluSrc1~0_combout\)) # (\Mux123~1_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001101110111001100110111011100110011001101110011001100110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(31),
	datab => \ALT_INV_Mux123~1_combout\,
	datac => \ALT_INV_R.curInst\(2),
	datad => \ALT_INV_vAluSrc1~0_combout\,
	dataf => \ALT_INV_R.curInst\(5),
	combout => \Mux123~3_combout\);

-- Location: FF_X61_Y5_N2
\RegFile[2][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(21),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][21]~q\);

-- Location: FF_X62_Y3_N50
\RegFile[5][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(21),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][21]~q\);

-- Location: MLABCELL_X59_Y5_N45
\RegFile[6][21]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[6][21]~feeder_combout\ = ( \R.regWriteData\(21) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(21),
	combout => \RegFile[6][21]~feeder_combout\);

-- Location: FF_X59_Y5_N46
\RegFile[6][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[6][21]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][21]~q\);

-- Location: LABCELL_X56_Y3_N39
\RegFile[4][21]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[4][21]~feeder_combout\ = ( \R.regWriteData\(21) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(21),
	combout => \RegFile[4][21]~feeder_combout\);

-- Location: FF_X56_Y3_N40
\RegFile[4][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[4][21]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][21]~q\);

-- Location: FF_X62_Y3_N19
\RegFile[7][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(21),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][21]~q\);

-- Location: LABCELL_X62_Y3_N18
\Mux69~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux69~0_combout\ = ( \RegFile[7][21]~q\ & ( \R.curInst\(15) & ( (\R.curInst\(16)) # (\RegFile[5][21]~q\) ) ) ) # ( !\RegFile[7][21]~q\ & ( \R.curInst\(15) & ( (\RegFile[5][21]~q\ & !\R.curInst\(16)) ) ) ) # ( \RegFile[7][21]~q\ & ( !\R.curInst\(15) & ( 
-- (!\R.curInst\(16) & ((\RegFile[4][21]~q\))) # (\R.curInst\(16) & (\RegFile[6][21]~q\)) ) ) ) # ( !\RegFile[7][21]~q\ & ( !\R.curInst\(15) & ( (!\R.curInst\(16) & ((\RegFile[4][21]~q\))) # (\R.curInst\(16) & (\RegFile[6][21]~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001111110011000000111111001101010000010100000101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[5][21]~q\,
	datab => \ALT_INV_RegFile[6][21]~q\,
	datac => \ALT_INV_R.curInst\(16),
	datad => \ALT_INV_RegFile[4][21]~q\,
	datae => \ALT_INV_RegFile[7][21]~q\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux69~0_combout\);

-- Location: LABCELL_X61_Y5_N18
\RegFile[1][21]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[1][21]~feeder_combout\ = ( \R.regWriteData\(21) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(21),
	combout => \RegFile[1][21]~feeder_combout\);

-- Location: FF_X61_Y5_N19
\RegFile[1][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[1][21]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][21]~q\);

-- Location: LABCELL_X62_Y3_N36
\Mux69~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux69~26_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (\R.curInst\(15) & (\RegFile[1][21]~q\))) # (\R.curInst\(17) & (((\Mux69~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & ((!\R.curInst\(15) & (((\RegFile[2][21]~q\)))) # 
-- (\R.curInst\(15) & (\RegFile[3][21]~q\)))) # (\R.curInst\(17) & ((((\Mux69~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000000000111010000000000000011111111110001110111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][21]~q\,
	datab => \ALT_INV_R.curInst\(15),
	datac => \ALT_INV_RegFile[2][21]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux69~0_combout\,
	datag => \ALT_INV_RegFile[1][21]~q\,
	combout => \Mux69~26_combout\);

-- Location: FF_X65_Y5_N2
\RegFile[13][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(21),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][21]~q\);

-- Location: MLABCELL_X65_Y5_N54
\RegFile[14][21]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[14][21]~feeder_combout\ = ( \R.regWriteData\(21) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(21),
	combout => \RegFile[14][21]~feeder_combout\);

-- Location: FF_X65_Y5_N56
\RegFile[14][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[14][21]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][21]~q\);

-- Location: FF_X65_Y5_N8
\RegFile[15][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(21),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][21]~q\);

-- Location: FF_X64_Y3_N38
\RegFile[9][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(21),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][21]~q\);

-- Location: FF_X64_Y3_N32
\RegFile[11][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(21),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][21]~q\);

-- Location: LABCELL_X64_Y3_N48
\RegFile[10][21]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[10][21]~feeder_combout\ = \R.regWriteData\(21)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110011001100110011001100110011001100110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.regWriteData\(21),
	combout => \RegFile[10][21]~feeder_combout\);

-- Location: FF_X64_Y3_N50
\RegFile[10][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[10][21]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][21]~q\);

-- Location: LABCELL_X56_Y3_N15
\RegFile[8][21]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[8][21]~feeder_combout\ = ( \R.regWriteData\(21) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(21),
	combout => \RegFile[8][21]~feeder_combout\);

-- Location: FF_X56_Y3_N16
\RegFile[8][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[8][21]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][21]~q\);

-- Location: LABCELL_X64_Y3_N30
\Mux69~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux69~14_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[8][21]~q\))) # (\R.curInst\(15) & (\RegFile[9][21]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[10][21]~q\))) # (\R.curInst\(15) & (\RegFile[11][21]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][21]~q\,
	datab => \ALT_INV_RegFile[11][21]~q\,
	datac => \ALT_INV_RegFile[10][21]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][21]~q\,
	combout => \Mux69~14_combout\);

-- Location: FF_X62_Y2_N46
\RegFile[12][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(21),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][21]~q\);

-- Location: MLABCELL_X65_Y5_N6
\Mux69~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux69~1_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux69~14_combout\))))) # (\R.curInst\(17) & (((!\Mux69~14_combout\ & ((\RegFile[12][21]~q\))) # (\Mux69~14_combout\ & (\RegFile[13][21]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux69~14_combout\)))) # (\R.curInst\(17) & ((!\Mux69~14_combout\ & (\RegFile[14][21]~q\)) # (\Mux69~14_combout\ & ((\RegFile[15][21]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][21]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[14][21]~q\,
	datad => \ALT_INV_RegFile[15][21]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux69~14_combout\,
	datag => \ALT_INV_RegFile[12][21]~q\,
	combout => \Mux69~1_combout\);

-- Location: FF_X66_Y3_N26
\RegFile[31][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(21),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][21]~q\);

-- Location: FF_X62_Y5_N32
\RegFile[29][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(21),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][21]~q\);

-- Location: FF_X66_Y3_N38
\RegFile[30][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(21),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][21]~q\);

-- Location: FF_X67_Y2_N2
\RegFile[27][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(21),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][21]~q\);

-- Location: FF_X67_Y2_N44
\RegFile[25][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(21),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][21]~q\);

-- Location: LABCELL_X67_Y2_N51
\RegFile[26][21]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[26][21]~feeder_combout\ = ( \R.regWriteData\(21) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(21),
	combout => \RegFile[26][21]~feeder_combout\);

-- Location: FF_X67_Y2_N53
\RegFile[26][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[26][21]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][21]~q\);

-- Location: LABCELL_X55_Y2_N27
\RegFile[24][21]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[24][21]~feeder_combout\ = ( \R.regWriteData\(21) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(21),
	combout => \RegFile[24][21]~feeder_combout\);

-- Location: FF_X55_Y2_N28
\RegFile[24][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[24][21]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][21]~q\);

-- Location: LABCELL_X67_Y2_N0
\Mux69~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux69~22_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[24][21]~q\))) # (\R.curInst\(15) & (\RegFile[25][21]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[26][21]~q\))) # (\R.curInst\(15) & (\RegFile[27][21]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[27][21]~q\,
	datab => \ALT_INV_RegFile[25][21]~q\,
	datac => \ALT_INV_RegFile[26][21]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][21]~q\,
	combout => \Mux69~22_combout\);

-- Location: LABCELL_X66_Y3_N18
\RegFile[28][21]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[28][21]~feeder_combout\ = \R.regWriteData\(21)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110011001100110011001100110011001100110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.regWriteData\(21),
	combout => \RegFile[28][21]~feeder_combout\);

-- Location: FF_X66_Y3_N19
\RegFile[28][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[28][21]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][21]~q\);

-- Location: LABCELL_X66_Y3_N24
\Mux69~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux69~9_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux69~22_combout\)))) # (\R.curInst\(17) & ((!\Mux69~22_combout\ & ((\RegFile[28][21]~q\))) # (\Mux69~22_combout\ & (\RegFile[29][21]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux69~22_combout\)))) # (\R.curInst\(17) & ((!\Mux69~22_combout\ & ((\RegFile[30][21]~q\))) # (\Mux69~22_combout\ & (\RegFile[31][21]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][21]~q\,
	datab => \ALT_INV_RegFile[29][21]~q\,
	datac => \ALT_INV_RegFile[30][21]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux69~22_combout\,
	datag => \ALT_INV_RegFile[28][21]~q\,
	combout => \Mux69~9_combout\);

-- Location: FF_X63_Y4_N50
\RegFile[23][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(21),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][21]~q\);

-- Location: FF_X59_Y1_N31
\RegFile[22][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(21),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][21]~q\);

-- Location: FF_X62_Y5_N14
\RegFile[21][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(21),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][21]~q\);

-- Location: FF_X63_Y4_N26
\RegFile[19][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(21),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][21]~q\);

-- Location: LABCELL_X63_Y5_N3
\RegFile[18][21]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[18][21]~feeder_combout\ = \R.regWriteData\(21)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101010101010101010101010101010101010101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.regWriteData\(21),
	combout => \RegFile[18][21]~feeder_combout\);

-- Location: FF_X63_Y5_N5
\RegFile[18][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][21]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][21]~q\);

-- Location: FF_X64_Y1_N14
\RegFile[17][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(21),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][21]~q\);

-- Location: LABCELL_X64_Y1_N0
\RegFile[16][21]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[16][21]~feeder_combout\ = ( \R.regWriteData\(21) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(21),
	combout => \RegFile[16][21]~feeder_combout\);

-- Location: FF_X64_Y1_N1
\RegFile[16][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[16][21]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][21]~q\);

-- Location: LABCELL_X63_Y4_N24
\Mux69~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux69~18_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & (\RegFile[16][21]~q\)) # (\R.curInst\(15) & ((\RegFile[17][21]~q\))))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & ((\RegFile[18][21]~q\))) # (\R.curInst\(15) & (\RegFile[19][21]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110000110011111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[19][21]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[18][21]~q\,
	datad => \ALT_INV_RegFile[17][21]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][21]~q\,
	combout => \Mux69~18_combout\);

-- Location: MLABCELL_X59_Y5_N15
\RegFile[20][21]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[20][21]~feeder_combout\ = ( \R.regWriteData\(21) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(21),
	combout => \RegFile[20][21]~feeder_combout\);

-- Location: FF_X59_Y5_N16
\RegFile[20][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[20][21]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][21]~q\);

-- Location: LABCELL_X63_Y4_N48
\Mux69~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux69~5_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux69~18_combout\)))) # (\R.curInst\(17) & ((!\Mux69~18_combout\ & (\RegFile[20][21]~q\)) # (\Mux69~18_combout\ & ((\RegFile[21][21]~q\)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) 
-- & ((((\Mux69~18_combout\))))) # (\R.curInst\(17) & (((!\Mux69~18_combout\ & ((\RegFile[22][21]~q\))) # (\Mux69~18_combout\ & (\RegFile[23][21]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111001100111111111101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[23][21]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[22][21]~q\,
	datad => \ALT_INV_RegFile[21][21]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux69~18_combout\,
	datag => \ALT_INV_RegFile[20][21]~q\,
	combout => \Mux69~5_combout\);

-- Location: MLABCELL_X65_Y5_N24
\Mux69~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux69~13_combout\ = ( \Mux69~9_combout\ & ( \Mux69~5_combout\ & ( ((!\R.curInst\(18) & (\Mux69~26_combout\)) # (\R.curInst\(18) & ((\Mux69~1_combout\)))) # (\R.curInst\(19)) ) ) ) # ( !\Mux69~9_combout\ & ( \Mux69~5_combout\ & ( (!\R.curInst\(19) & 
-- ((!\R.curInst\(18) & (\Mux69~26_combout\)) # (\R.curInst\(18) & ((\Mux69~1_combout\))))) # (\R.curInst\(19) & (!\R.curInst\(18))) ) ) ) # ( \Mux69~9_combout\ & ( !\Mux69~5_combout\ & ( (!\R.curInst\(19) & ((!\R.curInst\(18) & (\Mux69~26_combout\)) # 
-- (\R.curInst\(18) & ((\Mux69~1_combout\))))) # (\R.curInst\(19) & (\R.curInst\(18))) ) ) ) # ( !\Mux69~9_combout\ & ( !\Mux69~5_combout\ & ( (!\R.curInst\(19) & ((!\R.curInst\(18) & (\Mux69~26_combout\)) # (\R.curInst\(18) & ((\Mux69~1_combout\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000100000101010000110010011101101001100011011100101110101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(19),
	datab => \ALT_INV_R.curInst\(18),
	datac => \ALT_INV_Mux69~26_combout\,
	datad => \ALT_INV_Mux69~1_combout\,
	datae => \ALT_INV_Mux69~9_combout\,
	dataf => \ALT_INV_Mux69~5_combout\,
	combout => \Mux69~13_combout\);

-- Location: LABCELL_X74_Y5_N36
\Mux233~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux233~0_combout\ = ( \Mux69~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC[21]~DUPLICATE_q\))) ) ) # ( !\Mux69~13_combout\ & ( (!\vAluSrc1~1_combout\ & (\R.curPC[21]~DUPLICATE_q\ & \vAluSrc1~2_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000001100000000000000110011001100000011001100110000001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_vAluSrc1~1_combout\,
	datac => \ALT_INV_R.curPC[21]~DUPLICATE_q\,
	datad => \ALT_INV_vAluSrc1~2_combout\,
	dataf => \ALT_INV_Mux69~13_combout\,
	combout => \Mux233~0_combout\);

-- Location: FF_X72_Y5_N37
\R.aluData2[4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \NxR.aluData2[4]~20_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData2\(4));

-- Location: LABCELL_X77_Y5_N18
\Mux153~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux153~0_combout\ = ( \R.curInst\(8) & ( \R.curInst\(21) & ( ((\Mux53~0_combout\ & ((\Mux18~0_combout\) # (\Mux154~0_combout\)))) # (\Equal4~0_combout\) ) ) ) # ( !\R.curInst\(8) & ( \R.curInst\(21) & ( ((\Mux53~0_combout\ & \Mux154~0_combout\)) # 
-- (\Equal4~0_combout\) ) ) ) # ( \R.curInst\(8) & ( !\R.curInst\(21) & ( (\Mux53~0_combout\ & \Mux18~0_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000101010100011111000111110001111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux53~0_combout\,
	datab => \ALT_INV_Mux154~0_combout\,
	datac => \ALT_INV_Equal4~0_combout\,
	datad => \ALT_INV_Mux18~0_combout\,
	datae => \ALT_INV_R.curInst\(8),
	dataf => \ALT_INV_R.curInst\(21),
	combout => \Mux153~0_combout\);

-- Location: LABCELL_X80_Y2_N39
\Mux222~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux222~0_combout\ = ( !\R.curInst\(13) & ( \R.curInst\(12) ) ) # ( \R.curInst\(13) & ( !\R.curInst\(12) & ( !\R.curInst\(14) ) ) ) # ( !\R.curInst\(13) & ( !\R.curInst\(12) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111111100001111000011111111111111110000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.curInst\(14),
	datae => \ALT_INV_R.curInst\(13),
	dataf => \ALT_INV_R.curInst\(12),
	combout => \Mux222~0_combout\);

-- Location: IOIBUF_X89_Y21_N55
\avm_d_readdata[25]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(25),
	o => \avm_d_readdata[25]~input_o\);

-- Location: FF_X72_Y7_N10
\Add2~1_OTERM735_NEW_REG838\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux253~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Add2~1_OTERM735_OTERM839\);

-- Location: FF_X71_Y9_N26
\RegFile[31][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(0),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][0]~q\);

-- Location: FF_X70_Y9_N58
\RegFile[30][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(0),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][0]~q\);

-- Location: FF_X72_Y6_N44
\RegFile[29][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(0),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][0]~q\);

-- Location: FF_X67_Y4_N7
\RegFile[25][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(0),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][0]~q\);

-- Location: FF_X67_Y4_N52
\RegFile[26][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(0),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][0]~q\);

-- Location: FF_X67_Y4_N13
\RegFile[27][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(0),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][0]~q\);

-- Location: LABCELL_X55_Y6_N39
\RegFile[24][0]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[24][0]~feeder_combout\ = ( \R.regWriteData\(0) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(0),
	combout => \RegFile[24][0]~feeder_combout\);

-- Location: FF_X55_Y6_N40
\RegFile[24][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[24][0]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][0]~q\);

-- Location: LABCELL_X71_Y9_N9
\Mux90~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux90~22_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[24][0]~q\))) # (\R.curInst\(15) & (\RegFile[25][0]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & (\RegFile[26][0]~q\)) # (\R.curInst\(15) & ((\RegFile[27][0]~q\)))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001110111011101110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[25][0]~q\,
	datac => \ALT_INV_RegFile[26][0]~q\,
	datad => \ALT_INV_RegFile[27][0]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][0]~q\,
	combout => \Mux90~22_combout\);

-- Location: LABCELL_X71_Y8_N30
\RegFile[28][0]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[28][0]~feeder_combout\ = ( \R.regWriteData\(0) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(0),
	combout => \RegFile[28][0]~feeder_combout\);

-- Location: FF_X71_Y8_N31
\RegFile[28][0]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[28][0]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][0]~DUPLICATE_q\);

-- Location: LABCELL_X71_Y9_N24
\Mux90~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux90~9_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux90~22_combout\))))) # (\R.curInst\(17) & (((!\Mux90~22_combout\ & (\RegFile[28][0]~DUPLICATE_q\)) # (\Mux90~22_combout\ & ((\RegFile[29][0]~q\)))))) ) ) # ( \R.curInst\(16) & ( 
-- (!\R.curInst\(17) & ((((\Mux90~22_combout\))))) # (\R.curInst\(17) & (((!\Mux90~22_combout\ & ((\RegFile[30][0]~q\))) # (\Mux90~22_combout\ & (\RegFile[31][0]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110101010111111111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[31][0]~q\,
	datac => \ALT_INV_RegFile[30][0]~q\,
	datad => \ALT_INV_RegFile[29][0]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux90~22_combout\,
	datag => \ALT_INV_RegFile[28][0]~DUPLICATE_q\,
	combout => \Mux90~9_combout\);

-- Location: FF_X71_Y9_N50
\RegFile[2][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(0),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][0]~q\);

-- Location: LABCELL_X67_Y5_N27
\RegFile[4][0]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[4][0]~feeder_combout\ = ( \R.regWriteData\(0) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(0),
	combout => \RegFile[4][0]~feeder_combout\);

-- Location: FF_X67_Y5_N29
\RegFile[4][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[4][0]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][0]~q\);

-- Location: LABCELL_X67_Y6_N42
\RegFile[6][0]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[6][0]~feeder_combout\ = ( \R.regWriteData\(0) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(0),
	combout => \RegFile[6][0]~feeder_combout\);

-- Location: FF_X67_Y6_N43
\RegFile[6][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[6][0]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][0]~q\);

-- Location: LABCELL_X67_Y6_N12
\RegFile[5][0]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[5][0]~feeder_combout\ = ( \R.regWriteData\(0) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(0),
	combout => \RegFile[5][0]~feeder_combout\);

-- Location: FF_X67_Y6_N13
\RegFile[5][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[5][0]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][0]~q\);

-- Location: LABCELL_X67_Y6_N27
\RegFile[7][0]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[7][0]~feeder_combout\ = ( \R.regWriteData\(0) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(0),
	combout => \RegFile[7][0]~feeder_combout\);

-- Location: FF_X67_Y6_N28
\RegFile[7][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[7][0]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][0]~q\);

-- Location: LABCELL_X71_Y9_N57
\Mux90~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux90~0_combout\ = ( \R.curInst\(16) & ( \R.curInst\(15) & ( \RegFile[7][0]~q\ ) ) ) # ( !\R.curInst\(16) & ( \R.curInst\(15) & ( \RegFile[5][0]~q\ ) ) ) # ( \R.curInst\(16) & ( !\R.curInst\(15) & ( \RegFile[6][0]~q\ ) ) ) # ( !\R.curInst\(16) & ( 
-- !\R.curInst\(15) & ( \RegFile[4][0]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101001100110011001100001111000011110000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[4][0]~q\,
	datab => \ALT_INV_RegFile[6][0]~q\,
	datac => \ALT_INV_RegFile[5][0]~q\,
	datad => \ALT_INV_RegFile[7][0]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux90~0_combout\);

-- Location: LABCELL_X68_Y9_N3
\RegFile[1][0]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[1][0]~feeder_combout\ = ( \R.regWriteData\(0) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(0),
	combout => \RegFile[1][0]~feeder_combout\);

-- Location: FF_X68_Y9_N4
\RegFile[1][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[1][0]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][0]~q\);

-- Location: LABCELL_X71_Y9_N48
\Mux90~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux90~26_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((\RegFile[1][0]~q\ & ((\R.curInst\(15))))))) # (\R.curInst\(17) & ((((\Mux90~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[2][0]~q\))) # 
-- (\R.curInst\(15) & (\RegFile[3][0]~q\))))) # (\R.curInst\(17) & ((((\Mux90~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000001010101000010100101111100001010010111110010001001110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[3][0]~q\,
	datac => \ALT_INV_RegFile[2][0]~q\,
	datad => \ALT_INV_Mux90~0_combout\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[1][0]~q\,
	combout => \Mux90~26_combout\);

-- Location: FF_X70_Y8_N56
\RegFile[13][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(0),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][0]~q\);

-- Location: LABCELL_X56_Y8_N0
\RegFile[14][0]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[14][0]~feeder_combout\ = ( \R.regWriteData\(0) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(0),
	combout => \RegFile[14][0]~feeder_combout\);

-- Location: FF_X56_Y8_N1
\RegFile[14][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[14][0]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][0]~q\);

-- Location: FF_X66_Y8_N2
\RegFile[15][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(0),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][0]~q\);

-- Location: FF_X66_Y8_N14
\RegFile[11][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(0),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][0]~q\);

-- Location: LABCELL_X71_Y8_N36
\RegFile[9][0]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[9][0]~feeder_combout\ = ( \R.regWriteData\(0) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(0),
	combout => \RegFile[9][0]~feeder_combout\);

-- Location: FF_X71_Y8_N37
\RegFile[9][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[9][0]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][0]~q\);

-- Location: LABCELL_X64_Y8_N42
\RegFile[10][0]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[10][0]~feeder_combout\ = ( \R.regWriteData\(0) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(0),
	combout => \RegFile[10][0]~feeder_combout\);

-- Location: FF_X64_Y8_N43
\RegFile[10][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[10][0]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][0]~q\);

-- Location: LABCELL_X63_Y8_N54
\RegFile[8][0]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[8][0]~feeder_combout\ = ( \R.regWriteData\(0) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(0),
	combout => \RegFile[8][0]~feeder_combout\);

-- Location: FF_X63_Y8_N55
\RegFile[8][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[8][0]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][0]~q\);

-- Location: LABCELL_X70_Y8_N42
\Mux90~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux90~14_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[8][0]~q\))) # (\R.curInst\(15) & (\RegFile[9][0]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[10][0]~q\))) # (\R.curInst\(15) & (\RegFile[11][0]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[11][0]~q\,
	datab => \ALT_INV_RegFile[9][0]~q\,
	datac => \ALT_INV_RegFile[10][0]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][0]~q\,
	combout => \Mux90~14_combout\);

-- Location: FF_X70_Y8_N23
\RegFile[12][0]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(0),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][0]~DUPLICATE_q\);

-- Location: LABCELL_X70_Y8_N54
\Mux90~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux90~1_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux90~14_combout\))))) # (\R.curInst\(17) & (((!\Mux90~14_combout\ & ((\RegFile[12][0]~DUPLICATE_q\))) # (\Mux90~14_combout\ & (\RegFile[13][0]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- (!\R.curInst\(17) & ((((\Mux90~14_combout\))))) # (\R.curInst\(17) & (((!\Mux90~14_combout\ & (\RegFile[14][0]~q\)) # (\Mux90~14_combout\ & ((\RegFile[15][0]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110111011101110111010101011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[13][0]~q\,
	datac => \ALT_INV_RegFile[14][0]~q\,
	datad => \ALT_INV_RegFile[15][0]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux90~14_combout\,
	datag => \ALT_INV_RegFile[12][0]~DUPLICATE_q\,
	combout => \Mux90~1_combout\);

-- Location: FF_X70_Y5_N38
\RegFile[23][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(0),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][0]~q\);

-- Location: FF_X72_Y6_N2
\RegFile[21][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(0),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][0]~q\);

-- Location: FF_X74_Y4_N38
\RegFile[22][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(0),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][0]~q\);

-- Location: FF_X70_Y4_N1
\RegFile[19][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(0),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][0]~q\);

-- Location: LABCELL_X66_Y4_N15
\RegFile[18][0]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[18][0]~feeder_combout\ = ( \R.regWriteData\(0) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(0),
	combout => \RegFile[18][0]~feeder_combout\);

-- Location: FF_X66_Y4_N16
\RegFile[18][0]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][0]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][0]~DUPLICATE_q\);

-- Location: FF_X66_Y4_N50
\RegFile[17][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(0),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][0]~q\);

-- Location: FF_X74_Y4_N53
\RegFile[16][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(0),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][0]~q\);

-- Location: LABCELL_X70_Y4_N36
\Mux90~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux90~18_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & (\RegFile[16][0]~q\)) # (\R.curInst\(15) & ((\RegFile[17][0]~q\)))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & ((\RegFile[18][0]~DUPLICATE_q\))) # (\R.curInst\(15) & (\RegFile[19][0]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001010101111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[19][0]~q\,
	datac => \ALT_INV_RegFile[18][0]~DUPLICATE_q\,
	datad => \ALT_INV_RegFile[17][0]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][0]~q\,
	combout => \Mux90~18_combout\);

-- Location: FF_X75_Y4_N40
\RegFile[20][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(0),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][0]~q\);

-- Location: LABCELL_X70_Y5_N36
\Mux90~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux90~5_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux90~18_combout\)))) # (\R.curInst\(17) & ((!\Mux90~18_combout\ & ((\RegFile[20][0]~q\))) # (\Mux90~18_combout\ & (\RegFile[21][0]~q\))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) 
-- & (((\Mux90~18_combout\)))) # (\R.curInst\(17) & ((!\Mux90~18_combout\ & ((\RegFile[22][0]~q\))) # (\Mux90~18_combout\ & (\RegFile[23][0]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[23][0]~q\,
	datab => \ALT_INV_RegFile[21][0]~q\,
	datac => \ALT_INV_RegFile[22][0]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux90~18_combout\,
	datag => \ALT_INV_RegFile[20][0]~q\,
	combout => \Mux90~5_combout\);

-- Location: LABCELL_X71_Y9_N39
\Mux90~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux90~13_combout\ = ( \Mux90~1_combout\ & ( \Mux90~5_combout\ & ( (!\R.curInst\(19) & (((\Mux90~26_combout\) # (\R.curInst\(18))))) # (\R.curInst\(19) & (((!\R.curInst\(18))) # (\Mux90~9_combout\))) ) ) ) # ( !\Mux90~1_combout\ & ( \Mux90~5_combout\ & ( 
-- (!\R.curInst\(19) & (((!\R.curInst\(18) & \Mux90~26_combout\)))) # (\R.curInst\(19) & (((!\R.curInst\(18))) # (\Mux90~9_combout\))) ) ) ) # ( \Mux90~1_combout\ & ( !\Mux90~5_combout\ & ( (!\R.curInst\(19) & (((\Mux90~26_combout\) # (\R.curInst\(18))))) # 
-- (\R.curInst\(19) & (\Mux90~9_combout\ & (\R.curInst\(18)))) ) ) ) # ( !\Mux90~1_combout\ & ( !\Mux90~5_combout\ & ( (!\R.curInst\(19) & (((!\R.curInst\(18) & \Mux90~26_combout\)))) # (\R.curInst\(19) & (\Mux90~9_combout\ & (\R.curInst\(18)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000111000001000011011100110100110001111100010011110111111101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux90~9_combout\,
	datab => \ALT_INV_R.curInst\(19),
	datac => \ALT_INV_R.curInst\(18),
	datad => \ALT_INV_Mux90~26_combout\,
	datae => \ALT_INV_Mux90~1_combout\,
	dataf => \ALT_INV_Mux90~5_combout\,
	combout => \Mux90~13_combout\);

-- Location: MLABCELL_X72_Y7_N0
\Mux254~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux254~0_combout\ = ( \Mux90~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC[0]~DUPLICATE_q\))) ) ) # ( !\Mux90~13_combout\ & ( (!\vAluSrc1~1_combout\ & (\R.curPC[0]~DUPLICATE_q\ & \vAluSrc1~2_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000001100000000000000110011001100000011001100110000001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_vAluSrc1~1_combout\,
	datac => \ALT_INV_R.curPC[0]~DUPLICATE_q\,
	datad => \ALT_INV_vAluSrc1~2_combout\,
	dataf => \ALT_INV_Mux90~13_combout\,
	combout => \Mux254~0_combout\);

-- Location: FF_X72_Y7_N40
\Add2~1_OTERM735_NEW_REG836\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux254~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Add2~1_OTERM735_OTERM837\);

-- Location: MLABCELL_X78_Y6_N0
\Add1~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~2\ = CARRY(( \Add2~1_OTERM735_OTERM837\ ) + ( \R.aluData2\(0) ) + ( !VCC ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluData2\(0),
	datad => \ALT_INV_Add2~1_OTERM735_OTERM837\,
	cin => GND,
	cout => \Add1~2\);

-- Location: MLABCELL_X78_Y6_N3
\Add1~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~5_sumout\ = SUM(( \R.aluData2\(1) ) + ( \Add2~1_OTERM735_OTERM839\ ) + ( \Add1~2\ ))
-- \Add1~6\ = CARRY(( \R.aluData2\(1) ) + ( \Add2~1_OTERM735_OTERM839\ ) + ( \Add1~2\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Add2~1_OTERM735_OTERM839\,
	datad => \ALT_INV_R.aluData2\(1),
	cin => \Add1~2\,
	sumout => \Add1~5_sumout\,
	cout => \Add1~6\);

-- Location: LABCELL_X79_Y6_N0
\Add2~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~1_sumout\ = SUM(( !\R.aluData2\(0) $ (!\Add2~1_OTERM735_OTERM837\) ) + ( !VCC ) + ( !VCC ))
-- \Add2~2\ = CARRY(( !\R.aluData2\(0) $ (!\Add2~1_OTERM735_OTERM837\) ) + ( !VCC ) + ( !VCC ))
-- \Add2~3\ = SHARE((!\R.aluData2\(0)) # (\Add2~1_OTERM735_OTERM837\))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111111100000000000000000000111111110000",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluData2\(0),
	datad => \ALT_INV_Add2~1_OTERM735_OTERM837\,
	cin => GND,
	sharein => GND,
	sumout => \Add2~1_sumout\,
	cout => \Add2~2\,
	shareout => \Add2~3\);

-- Location: LABCELL_X79_Y6_N3
\Add2~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~5_sumout\ = SUM(( !\Add2~1_OTERM735_OTERM839\ $ (\R.aluData2\(1)) ) + ( \Add2~3\ ) + ( \Add2~2\ ))
-- \Add2~6\ = CARRY(( !\Add2~1_OTERM735_OTERM839\ $ (\R.aluData2\(1)) ) + ( \Add2~3\ ) + ( \Add2~2\ ))
-- \Add2~7\ = SHARE((\Add2~1_OTERM735_OTERM839\ & !\R.aluData2\(1)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000000000000000000000001111000000001111",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Add2~1_OTERM735_OTERM839\,
	datad => \ALT_INV_R.aluData2\(1),
	cin => \Add2~2\,
	sharein => \Add2~3\,
	sumout => \Add2~5_sumout\,
	cout => \Add2~6\,
	shareout => \Add2~7\);

-- Location: LABCELL_X77_Y5_N0
\Mux151~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux151~0_combout\ = ( \R.curInst\(23) & ( \R.curInst\(10) & ( ((\Mux53~0_combout\ & ((\Mux18~0_combout\) # (\Mux154~0_combout\)))) # (\Equal4~0_combout\) ) ) ) # ( !\R.curInst\(23) & ( \R.curInst\(10) & ( (\Mux53~0_combout\ & \Mux18~0_combout\) ) ) ) # ( 
-- \R.curInst\(23) & ( !\R.curInst\(10) & ( ((\Mux53~0_combout\ & \Mux154~0_combout\)) # (\Equal4~0_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000111110001111100000000010101010001111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux53~0_combout\,
	datab => \ALT_INV_Mux154~0_combout\,
	datac => \ALT_INV_Equal4~0_combout\,
	datad => \ALT_INV_Mux18~0_combout\,
	datae => \ALT_INV_R.curInst\(23),
	dataf => \ALT_INV_R.curInst\(10),
	combout => \Mux151~0_combout\);

-- Location: FF_X70_Y7_N41
\RegFile[21][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(3),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][3]~q\);

-- Location: FF_X71_Y5_N50
\RegFile[23][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(3),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][3]~q\);

-- Location: LABCELL_X63_Y9_N39
\RegFile[22][3]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[22][3]~feeder_combout\ = ( \R.regWriteData\(3) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(3),
	combout => \RegFile[22][3]~feeder_combout\);

-- Location: FF_X63_Y9_N40
\RegFile[22][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[22][3]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][3]~q\);

-- Location: FF_X70_Y4_N38
\RegFile[17][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(3),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][3]~q\);

-- Location: FF_X66_Y4_N31
\RegFile[18][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(3),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][3]~q\);

-- Location: LABCELL_X70_Y4_N57
\RegFile[19][3]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[19][3]~feeder_combout\ = ( \R.regWriteData\(3) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(3),
	combout => \RegFile[19][3]~feeder_combout\);

-- Location: FF_X70_Y4_N58
\RegFile[19][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[19][3]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][3]~q\);

-- Location: LABCELL_X68_Y9_N9
\RegFile[16][3]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[16][3]~feeder_combout\ = ( \R.regWriteData\(3) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(3),
	combout => \RegFile[16][3]~feeder_combout\);

-- Location: FF_X68_Y9_N10
\RegFile[16][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[16][3]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][3]~q\);

-- Location: LABCELL_X70_Y7_N30
\Mux87~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux87~18_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[16][3]~q\))) # (\R.curInst\(15) & (\RegFile[17][3]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & (\RegFile[18][3]~q\)) # (\R.curInst\(15) & ((\RegFile[19][3]~q\))))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[17][3]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[18][3]~q\,
	datad => \ALT_INV_RegFile[19][3]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][3]~q\,
	combout => \Mux87~18_combout\);

-- Location: FF_X68_Y6_N38
\RegFile[20][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(3),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][3]~q\);

-- Location: LABCELL_X71_Y5_N48
\Mux87~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux87~5_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux87~18_combout\)))) # (\R.curInst\(17) & ((!\Mux87~18_combout\ & ((\RegFile[20][3]~q\))) # (\Mux87~18_combout\ & (\RegFile[21][3]~q\))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) 
-- & (((\Mux87~18_combout\)))) # (\R.curInst\(17) & ((!\Mux87~18_combout\ & ((\RegFile[22][3]~q\))) # (\Mux87~18_combout\ & (\RegFile[23][3]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][3]~q\,
	datab => \ALT_INV_RegFile[23][3]~q\,
	datac => \ALT_INV_RegFile[22][3]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux87~18_combout\,
	datag => \ALT_INV_RegFile[20][3]~q\,
	combout => \Mux87~5_combout\);

-- Location: FF_X70_Y7_N26
\RegFile[3][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(3),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][3]~q\);

-- Location: FF_X71_Y5_N44
\RegFile[2][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(3),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][3]~q\);

-- Location: LABCELL_X60_Y4_N30
\RegFile[4][3]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[4][3]~feeder_combout\ = ( \R.regWriteData\(3) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(3),
	combout => \RegFile[4][3]~feeder_combout\);

-- Location: FF_X60_Y4_N31
\RegFile[4][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[4][3]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][3]~q\);

-- Location: MLABCELL_X65_Y7_N27
\RegFile[5][3]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[5][3]~feeder_combout\ = ( \R.regWriteData\(3) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(3),
	combout => \RegFile[5][3]~feeder_combout\);

-- Location: FF_X65_Y7_N29
\RegFile[5][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[5][3]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][3]~q\);

-- Location: FF_X68_Y4_N44
\RegFile[6][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(3),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][3]~q\);

-- Location: FF_X68_Y4_N50
\RegFile[7][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(3),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][3]~q\);

-- Location: LABCELL_X68_Y4_N48
\Mux87~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux87~0_combout\ = ( \RegFile[7][3]~q\ & ( \R.curInst\(15) & ( (\RegFile[5][3]~q\) # (\R.curInst\(16)) ) ) ) # ( !\RegFile[7][3]~q\ & ( \R.curInst\(15) & ( (!\R.curInst\(16) & \RegFile[5][3]~q\) ) ) ) # ( \RegFile[7][3]~q\ & ( !\R.curInst\(15) & ( 
-- (!\R.curInst\(16) & (\RegFile[4][3]~q\)) # (\R.curInst\(16) & ((\RegFile[6][3]~q\))) ) ) ) # ( !\RegFile[7][3]~q\ & ( !\R.curInst\(15) & ( (!\R.curInst\(16) & (\RegFile[4][3]~q\)) # (\R.curInst\(16) & ((\RegFile[6][3]~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100010001110111010001000111011100001100000011000011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[4][3]~q\,
	datab => \ALT_INV_R.curInst\(16),
	datac => \ALT_INV_RegFile[5][3]~q\,
	datad => \ALT_INV_RegFile[6][3]~q\,
	datae => \ALT_INV_RegFile[7][3]~q\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux87~0_combout\);

-- Location: LABCELL_X68_Y9_N51
\RegFile[1][3]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[1][3]~feeder_combout\ = ( \R.regWriteData\(3) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(3),
	combout => \RegFile[1][3]~feeder_combout\);

-- Location: FF_X68_Y9_N52
\RegFile[1][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[1][3]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][3]~q\);

-- Location: LABCELL_X71_Y5_N42
\Mux87~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux87~26_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (\R.curInst\(15) & (\RegFile[1][3]~q\))) # (\R.curInst\(17) & (((\Mux87~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & ((!\R.curInst\(15) & (((\RegFile[2][3]~q\)))) # 
-- (\R.curInst\(15) & (\RegFile[3][3]~q\)))) # (\R.curInst\(17) & ((((\Mux87~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000000000110110000000000000101111111110001101111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(15),
	datab => \ALT_INV_RegFile[3][3]~q\,
	datac => \ALT_INV_RegFile[2][3]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux87~0_combout\,
	datag => \ALT_INV_RegFile[1][3]~q\,
	combout => \Mux87~26_combout\);

-- Location: FF_X66_Y1_N41
\RegFile[15][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(3),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][3]~q\);

-- Location: LABCELL_X66_Y1_N54
\RegFile[14][3]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[14][3]~feeder_combout\ = ( \R.regWriteData\(3) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(3),
	combout => \RegFile[14][3]~feeder_combout\);

-- Location: FF_X66_Y1_N55
\RegFile[14][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[14][3]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][3]~q\);

-- Location: FF_X65_Y1_N20
\RegFile[11][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(3),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][3]~q\);

-- Location: FF_X66_Y1_N26
\RegFile[9][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(3),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][3]~q\);

-- Location: FF_X57_Y1_N37
\RegFile[10][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(3),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][3]~q\);

-- Location: FF_X66_Y5_N28
\RegFile[8][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(3),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][3]~q\);

-- Location: MLABCELL_X65_Y1_N18
\Mux87~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux87~14_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[8][3]~q\))) # (\R.curInst\(15) & (\RegFile[9][3]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[10][3]~q\))) # (\R.curInst\(15) & (\RegFile[11][3]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[11][3]~q\,
	datab => \ALT_INV_RegFile[9][3]~q\,
	datac => \ALT_INV_RegFile[10][3]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][3]~q\,
	combout => \Mux87~14_combout\);

-- Location: FF_X57_Y1_N52
\RegFile[12][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(3),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][3]~q\);

-- Location: MLABCELL_X65_Y1_N30
\Mux87~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux87~1_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux87~14_combout\)))) # (\R.curInst\(17) & ((!\Mux87~14_combout\ & ((\RegFile[12][3]~q\))) # (\Mux87~14_combout\ & (\RegFile[13][3]~q\))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) 
-- & (((\Mux87~14_combout\)))) # (\R.curInst\(17) & ((!\Mux87~14_combout\ & ((\RegFile[14][3]~q\))) # (\Mux87~14_combout\ & (\RegFile[15][3]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][3]~q\,
	datab => \ALT_INV_RegFile[13][3]~q\,
	datac => \ALT_INV_RegFile[14][3]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux87~14_combout\,
	datag => \ALT_INV_RegFile[12][3]~q\,
	combout => \Mux87~1_combout\);

-- Location: FF_X68_Y6_N14
\RegFile[29][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(3),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][3]~q\);

-- Location: FF_X65_Y4_N8
\RegFile[31][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(3),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][3]~q\);

-- Location: FF_X60_Y6_N22
\RegFile[30][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(3),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][3]~q\);

-- Location: FF_X65_Y4_N44
\RegFile[25][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(3),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][3]~q\);

-- Location: FF_X67_Y4_N59
\RegFile[26][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(3),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][3]~q\);

-- Location: FF_X65_Y4_N32
\RegFile[27][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(3),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][3]~q\);

-- Location: LABCELL_X60_Y4_N6
\RegFile[24][3]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[24][3]~feeder_combout\ = ( \R.regWriteData\(3) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(3),
	combout => \RegFile[24][3]~feeder_combout\);

-- Location: FF_X60_Y4_N7
\RegFile[24][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[24][3]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][3]~q\);

-- Location: MLABCELL_X65_Y4_N30
\Mux87~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux87~22_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[24][3]~q\))) # (\R.curInst\(15) & (\RegFile[25][3]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & (\RegFile[26][3]~q\)) # (\R.curInst\(15) & ((\RegFile[27][3]~q\)))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001110111011101110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[25][3]~q\,
	datac => \ALT_INV_RegFile[26][3]~q\,
	datad => \ALT_INV_RegFile[27][3]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][3]~q\,
	combout => \Mux87~22_combout\);

-- Location: MLABCELL_X65_Y9_N57
\RegFile[28][3]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[28][3]~feeder_combout\ = ( \R.regWriteData\(3) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(3),
	combout => \RegFile[28][3]~feeder_combout\);

-- Location: FF_X65_Y9_N59
\RegFile[28][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[28][3]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][3]~q\);

-- Location: MLABCELL_X65_Y4_N6
\Mux87~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux87~9_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux87~22_combout\)))) # (\R.curInst\(17) & ((!\Mux87~22_combout\ & ((\RegFile[28][3]~q\))) # (\Mux87~22_combout\ & (\RegFile[29][3]~q\))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) 
-- & (((\Mux87~22_combout\)))) # (\R.curInst\(17) & ((!\Mux87~22_combout\ & ((\RegFile[30][3]~q\))) # (\Mux87~22_combout\ & (\RegFile[31][3]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[29][3]~q\,
	datab => \ALT_INV_RegFile[31][3]~q\,
	datac => \ALT_INV_RegFile[30][3]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux87~22_combout\,
	datag => \ALT_INV_RegFile[28][3]~q\,
	combout => \Mux87~9_combout\);

-- Location: LABCELL_X71_Y5_N24
\Mux87~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux87~13_combout\ = ( \Mux87~1_combout\ & ( \Mux87~9_combout\ & ( ((!\R.curInst\(19) & ((\Mux87~26_combout\))) # (\R.curInst\(19) & (\Mux87~5_combout\))) # (\R.curInst\(18)) ) ) ) # ( !\Mux87~1_combout\ & ( \Mux87~9_combout\ & ( (!\R.curInst\(19) & 
-- (((\Mux87~26_combout\ & !\R.curInst\(18))))) # (\R.curInst\(19) & (((\R.curInst\(18))) # (\Mux87~5_combout\))) ) ) ) # ( \Mux87~1_combout\ & ( !\Mux87~9_combout\ & ( (!\R.curInst\(19) & (((\R.curInst\(18)) # (\Mux87~26_combout\)))) # (\R.curInst\(19) & 
-- (\Mux87~5_combout\ & ((!\R.curInst\(18))))) ) ) ) # ( !\Mux87~1_combout\ & ( !\Mux87~9_combout\ & ( (!\R.curInst\(18) & ((!\R.curInst\(19) & ((\Mux87~26_combout\))) # (\R.curInst\(19) & (\Mux87~5_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011010100000000001101011111000000110101000011110011010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux87~5_combout\,
	datab => \ALT_INV_Mux87~26_combout\,
	datac => \ALT_INV_R.curInst\(19),
	datad => \ALT_INV_R.curInst\(18),
	datae => \ALT_INV_Mux87~1_combout\,
	dataf => \ALT_INV_Mux87~9_combout\,
	combout => \Mux87~13_combout\);

-- Location: MLABCELL_X72_Y7_N54
\Mux251~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux251~0_combout\ = ( \Mux87~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC\(3)))) ) ) # ( !\Mux87~13_combout\ & ( (\R.curPC\(3) & (!\vAluSrc1~1_combout\ & \vAluSrc1~2_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110000000000000011000011110000001100001111000000110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.curPC\(3),
	datac => \ALT_INV_vAluSrc1~1_combout\,
	datad => \ALT_INV_vAluSrc1~2_combout\,
	dataf => \ALT_INV_Mux87~13_combout\,
	combout => \Mux251~0_combout\);

-- Location: FF_X71_Y7_N38
\RegFile[13][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(2),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][2]~q\);

-- Location: FF_X66_Y10_N7
\RegFile[14][2]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(2),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][2]~DUPLICATE_q\);

-- Location: FF_X72_Y8_N20
\RegFile[15][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(2),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][2]~q\);

-- Location: LABCELL_X66_Y8_N54
\RegFile[11][2]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[11][2]~feeder_combout\ = ( \R.regWriteData\(2) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(2),
	combout => \RegFile[11][2]~feeder_combout\);

-- Location: FF_X66_Y8_N55
\RegFile[11][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[11][2]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][2]~q\);

-- Location: LABCELL_X56_Y8_N39
\RegFile[10][2]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[10][2]~feeder_combout\ = ( \R.regWriteData\(2) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(2),
	combout => \RegFile[10][2]~feeder_combout\);

-- Location: FF_X56_Y8_N40
\RegFile[10][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[10][2]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][2]~q\);

-- Location: LABCELL_X66_Y8_N48
\RegFile[9][2]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[9][2]~feeder_combout\ = ( \R.regWriteData\(2) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(2),
	combout => \RegFile[9][2]~feeder_combout\);

-- Location: FF_X66_Y8_N49
\RegFile[9][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[9][2]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][2]~q\);

-- Location: LABCELL_X63_Y8_N42
\RegFile[8][2]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[8][2]~feeder_combout\ = ( \R.regWriteData\(2) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(2),
	combout => \RegFile[8][2]~feeder_combout\);

-- Location: FF_X63_Y8_N43
\RegFile[8][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[8][2]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][2]~q\);

-- Location: MLABCELL_X72_Y8_N33
\Mux88~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux88~14_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & (\RegFile[8][2]~q\)) # (\R.curInst\(15) & ((\RegFile[9][2]~q\))))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & ((\RegFile[10][2]~q\))) # (\R.curInst\(15) & (\RegFile[11][2]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110000110011111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[11][2]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[10][2]~q\,
	datad => \ALT_INV_RegFile[9][2]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][2]~q\,
	combout => \Mux88~14_combout\);

-- Location: FF_X66_Y10_N4
\RegFile[12][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(2),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][2]~q\);

-- Location: MLABCELL_X72_Y8_N18
\Mux88~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux88~1_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux88~14_combout\))))) # (\R.curInst\(17) & (((!\Mux88~14_combout\ & ((\RegFile[12][2]~q\))) # (\Mux88~14_combout\ & (\RegFile[13][2]~q\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) 
-- & ((((\Mux88~14_combout\))))) # (\R.curInst\(17) & (((!\Mux88~14_combout\ & (\RegFile[14][2]~DUPLICATE_q\)) # (\Mux88~14_combout\ & ((\RegFile[15][2]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110111011101110111010101011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[13][2]~q\,
	datac => \ALT_INV_RegFile[14][2]~DUPLICATE_q\,
	datad => \ALT_INV_RegFile[15][2]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux88~14_combout\,
	datag => \ALT_INV_RegFile[12][2]~q\,
	combout => \Mux88~1_combout\);

-- Location: FF_X68_Y8_N50
\RegFile[31][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(2),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][2]~q\);

-- Location: FF_X70_Y10_N53
\RegFile[29][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(2),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][2]~q\);

-- Location: FF_X66_Y10_N37
\RegFile[30][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(2),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][2]~q\);

-- Location: FF_X67_Y10_N37
\RegFile[27][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(2),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][2]~q\);

-- Location: FF_X70_Y10_N44
\RegFile[25][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(2),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][2]~q\);

-- Location: FF_X63_Y9_N16
\RegFile[26][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(2),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][2]~q\);

-- Location: LABCELL_X64_Y6_N57
\RegFile[24][2]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[24][2]~feeder_combout\ = \R.regWriteData\(2)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101010101010101010101010101010101010101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.regWriteData\(2),
	combout => \RegFile[24][2]~feeder_combout\);

-- Location: FF_X64_Y6_N58
\RegFile[24][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[24][2]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][2]~q\);

-- Location: LABCELL_X68_Y8_N42
\Mux88~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux88~22_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[24][2]~q\))) # (\R.curInst\(15) & (\RegFile[25][2]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[26][2]~q\))) # (\R.curInst\(15) & (\RegFile[27][2]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[27][2]~q\,
	datab => \ALT_INV_RegFile[25][2]~q\,
	datac => \ALT_INV_RegFile[26][2]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][2]~q\,
	combout => \Mux88~22_combout\);

-- Location: LABCELL_X70_Y9_N18
\RegFile[28][2]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[28][2]~feeder_combout\ = ( \R.regWriteData\(2) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(2),
	combout => \RegFile[28][2]~feeder_combout\);

-- Location: FF_X70_Y9_N19
\RegFile[28][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[28][2]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][2]~q\);

-- Location: LABCELL_X68_Y8_N48
\Mux88~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux88~9_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux88~22_combout\)))) # (\R.curInst\(17) & ((!\Mux88~22_combout\ & ((\RegFile[28][2]~q\))) # (\Mux88~22_combout\ & (\RegFile[29][2]~q\))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) 
-- & (((\Mux88~22_combout\)))) # (\R.curInst\(17) & ((!\Mux88~22_combout\ & ((\RegFile[30][2]~q\))) # (\Mux88~22_combout\ & (\RegFile[31][2]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][2]~q\,
	datab => \ALT_INV_RegFile[29][2]~q\,
	datac => \ALT_INV_RegFile[30][2]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux88~22_combout\,
	datag => \ALT_INV_RegFile[28][2]~q\,
	combout => \Mux88~9_combout\);

-- Location: FF_X72_Y8_N2
\RegFile[21][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(2),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][2]~q\);

-- Location: FF_X72_Y8_N29
\RegFile[23][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(2),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][2]~q\);

-- Location: FF_X73_Y10_N43
\RegFile[22][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(2),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][2]~q\);

-- Location: MLABCELL_X65_Y8_N54
\RegFile[17][2]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[17][2]~feeder_combout\ = ( \R.regWriteData\(2) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(2),
	combout => \RegFile[17][2]~feeder_combout\);

-- Location: FF_X65_Y8_N55
\RegFile[17][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[17][2]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][2]~q\);

-- Location: LABCELL_X64_Y10_N21
\RegFile[18][2]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[18][2]~feeder_combout\ = ( \R.regWriteData\(2) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(2),
	combout => \RegFile[18][2]~feeder_combout\);

-- Location: FF_X64_Y10_N22
\RegFile[18][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][2]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][2]~q\);

-- Location: MLABCELL_X65_Y8_N48
\RegFile[19][2]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[19][2]~feeder_combout\ = ( \R.regWriteData\(2) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(2),
	combout => \RegFile[19][2]~feeder_combout\);

-- Location: FF_X65_Y8_N49
\RegFile[19][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[19][2]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][2]~q\);

-- Location: FF_X63_Y9_N31
\RegFile[16][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(2),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][2]~q\);

-- Location: MLABCELL_X72_Y8_N12
\Mux88~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux88~18_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[16][2]~q\))) # (\R.curInst\(15) & (\RegFile[17][2]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & (\RegFile[18][2]~q\)) # (\R.curInst\(15) & ((\RegFile[19][2]~q\)))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001110111011101110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[17][2]~q\,
	datac => \ALT_INV_RegFile[18][2]~q\,
	datad => \ALT_INV_RegFile[19][2]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][2]~q\,
	combout => \Mux88~18_combout\);

-- Location: FF_X73_Y10_N40
\RegFile[20][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(2),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][2]~q\);

-- Location: MLABCELL_X72_Y8_N27
\Mux88~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux88~5_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux88~18_combout\)))) # (\R.curInst\(17) & ((!\Mux88~18_combout\ & ((\RegFile[20][2]~q\))) # (\Mux88~18_combout\ & (\RegFile[21][2]~q\))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) 
-- & (((\Mux88~18_combout\)))) # (\R.curInst\(17) & ((!\Mux88~18_combout\ & ((\RegFile[22][2]~q\))) # (\Mux88~18_combout\ & (\RegFile[23][2]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][2]~q\,
	datab => \ALT_INV_RegFile[23][2]~q\,
	datac => \ALT_INV_RegFile[22][2]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux88~18_combout\,
	datag => \ALT_INV_RegFile[20][2]~q\,
	combout => \Mux88~5_combout\);

-- Location: FF_X66_Y9_N56
\RegFile[6][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(2),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][2]~q\);

-- Location: FF_X57_Y7_N49
\RegFile[4][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(2),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][2]~q\);

-- Location: LABCELL_X62_Y9_N15
\RegFile[5][2]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[5][2]~feeder_combout\ = ( \R.regWriteData\(2) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(2),
	combout => \RegFile[5][2]~feeder_combout\);

-- Location: FF_X62_Y9_N16
\RegFile[5][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[5][2]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][2]~q\);

-- Location: FF_X66_Y9_N49
\RegFile[7][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(2),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][2]~q\);

-- Location: LABCELL_X66_Y9_N48
\Mux88~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux88~0_combout\ = ( \RegFile[7][2]~q\ & ( \R.curInst\(15) & ( (\RegFile[5][2]~q\) # (\R.curInst\(16)) ) ) ) # ( !\RegFile[7][2]~q\ & ( \R.curInst\(15) & ( (!\R.curInst\(16) & \RegFile[5][2]~q\) ) ) ) # ( \RegFile[7][2]~q\ & ( !\R.curInst\(15) & ( 
-- (!\R.curInst\(16) & ((\RegFile[4][2]~q\))) # (\R.curInst\(16) & (\RegFile[6][2]~q\)) ) ) ) # ( !\RegFile[7][2]~q\ & ( !\R.curInst\(15) & ( (!\R.curInst\(16) & ((\RegFile[4][2]~q\))) # (\R.curInst\(16) & (\RegFile[6][2]~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011010100110101001101010011010100000000111100000000111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[6][2]~q\,
	datab => \ALT_INV_RegFile[4][2]~q\,
	datac => \ALT_INV_R.curInst\(16),
	datad => \ALT_INV_RegFile[5][2]~q\,
	datae => \ALT_INV_RegFile[7][2]~q\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux88~0_combout\);

-- Location: FF_X71_Y7_N8
\RegFile[3][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(2),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][2]~q\);

-- Location: LABCELL_X64_Y10_N51
\RegFile[1][2]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[1][2]~feeder_combout\ = ( \R.regWriteData\(2) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(2),
	combout => \RegFile[1][2]~feeder_combout\);

-- Location: FF_X64_Y10_N52
\RegFile[1][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[1][2]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][2]~q\);

-- Location: LABCELL_X66_Y9_N0
\Mux88~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux88~26_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\RegFile[1][2]~q\ & \R.curInst\(15))))) # (\R.curInst\(17) & (\Mux88~0_combout\))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[2][2]~q\))) # 
-- (\R.curInst\(15) & (\RegFile[3][2]~q\))))) # (\R.curInst\(17) & (\Mux88~0_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000001010101000011110101010100001111010101010011001101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux88~0_combout\,
	datab => \ALT_INV_RegFile[3][2]~q\,
	datac => \ALT_INV_RegFile[2][2]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[1][2]~q\,
	combout => \Mux88~26_combout\);

-- Location: MLABCELL_X72_Y8_N39
\Mux88~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux88~13_combout\ = ( \Mux88~5_combout\ & ( \Mux88~26_combout\ & ( (!\R.curInst\(18)) # ((!\R.curInst\(19) & (\Mux88~1_combout\)) # (\R.curInst\(19) & ((\Mux88~9_combout\)))) ) ) ) # ( !\Mux88~5_combout\ & ( \Mux88~26_combout\ & ( (!\R.curInst\(19) & 
-- (((!\R.curInst\(18))) # (\Mux88~1_combout\))) # (\R.curInst\(19) & (((\Mux88~9_combout\ & \R.curInst\(18))))) ) ) ) # ( \Mux88~5_combout\ & ( !\Mux88~26_combout\ & ( (!\R.curInst\(19) & (\Mux88~1_combout\ & ((\R.curInst\(18))))) # (\R.curInst\(19) & 
-- (((!\R.curInst\(18)) # (\Mux88~9_combout\)))) ) ) ) # ( !\Mux88~5_combout\ & ( !\Mux88~26_combout\ & ( (\R.curInst\(18) & ((!\R.curInst\(19) & (\Mux88~1_combout\)) # (\R.curInst\(19) & ((\Mux88~9_combout\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001000111001100110100011111001100010001111111111101000111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux88~1_combout\,
	datab => \ALT_INV_R.curInst\(19),
	datac => \ALT_INV_Mux88~9_combout\,
	datad => \ALT_INV_R.curInst\(18),
	datae => \ALT_INV_Mux88~5_combout\,
	dataf => \ALT_INV_Mux88~26_combout\,
	combout => \Mux88~13_combout\);

-- Location: MLABCELL_X72_Y7_N15
\Mux252~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux252~0_combout\ = ( \Mux88~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC\(2)))) ) ) # ( !\Mux88~13_combout\ & ( (\vAluSrc1~2_combout\ & (!\vAluSrc1~1_combout\ & \R.curPC\(2))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110000000000000011000011000000111100001100000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_vAluSrc1~2_combout\,
	datac => \ALT_INV_vAluSrc1~1_combout\,
	datad => \ALT_INV_R.curPC\(2),
	dataf => \ALT_INV_Mux88~13_combout\,
	combout => \Mux252~0_combout\);

-- Location: MLABCELL_X72_Y7_N48
\ShiftLeft0~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~3_combout\ = ( \NxR.aluData2[0]~16_combout\ & ( \Mux252~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\) # (\Mux254~0_combout\) ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( \Mux252~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & 
-- ((\Mux251~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux253~0_combout\)) ) ) ) # ( \NxR.aluData2[0]~16_combout\ & ( !\Mux252~0_combout\ & ( (\NxR.aluData2[1]~17_combout\ & \Mux254~0_combout\) ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( 
-- !\Mux252~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((\Mux251~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux253~0_combout\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000111011101000000110000001100010001110111011100111111001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux253~0_combout\,
	datab => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datac => \ALT_INV_Mux254~0_combout\,
	datad => \ALT_INV_Mux251~0_combout\,
	datae => \ALT_INV_NxR.aluData2[0]~16_combout\,
	dataf => \ALT_INV_Mux252~0_combout\,
	combout => \ShiftLeft0~3_combout\);

-- Location: FF_X72_Y7_N49
\ShiftLeft0~3_NEW_REG222\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~3_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~3_OTERM223\);

-- Location: FF_X73_Y6_N28
\R.aluOp.ALUOpXor~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.aluOp.ALUOpXor_OTERM355\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluOp.ALUOpXor~DUPLICATE_q\);

-- Location: LABCELL_X77_Y6_N9
\Mux23~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux23~0_combout\ = ( \R.curInst\(13) & ( (\R.aluOp.ALUOpXor~DUPLICATE_q\ & \R.curInst\(6)) ) ) # ( !\R.curInst\(13) & ( (!\R.aluOp.ALUOpXor~DUPLICATE_q\ & (!\R.curInst\(12) & ((\Mux21~0_combout\)))) # (\R.aluOp.ALUOpXor~DUPLICATE_q\ & (((!\R.curInst\(12) 
-- & \Mux21~0_combout\)) # (\R.curInst\(6)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010111001101000001011100110100000101000001010000010100000101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpXor~DUPLICATE_q\,
	datab => \ALT_INV_R.curInst\(12),
	datac => \ALT_INV_R.curInst\(6),
	datad => \ALT_INV_Mux21~0_combout\,
	dataf => \ALT_INV_R.curInst\(13),
	combout => \Mux23~0_combout\);

-- Location: LABCELL_X77_Y6_N48
\Mux23~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux23~1_combout\ = ( \R.aluOp.ALUOpXor~DUPLICATE_q\ & ( \Mux23~0_combout\ & ( ((!\R.curInst\(3) & (!\Mux26~0_combout\)) # (\R.curInst\(3) & ((!\Mux123~0_combout\)))) # (\R.curInst\(4)) ) ) ) # ( !\R.aluOp.ALUOpXor~DUPLICATE_q\ & ( \Mux23~0_combout\ & ( 
-- (\R.curInst\(4) & !\R.curInst\(3)) ) ) ) # ( \R.aluOp.ALUOpXor~DUPLICATE_q\ & ( !\Mux23~0_combout\ & ( (!\R.curInst\(4) & ((!\R.curInst\(3) & (!\Mux26~0_combout\)) # (\R.curInst\(3) & ((!\Mux123~0_combout\))))) # (\R.curInst\(4) & (((\R.curInst\(3))))) ) 
-- ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000100011111000010101010000010100001101111111010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(4),
	datab => \ALT_INV_Mux26~0_combout\,
	datac => \ALT_INV_R.curInst\(3),
	datad => \ALT_INV_Mux123~0_combout\,
	datae => \ALT_INV_R.aluOp.ALUOpXor~DUPLICATE_q\,
	dataf => \ALT_INV_Mux23~0_combout\,
	combout => \Mux23~1_combout\);

-- Location: FF_X73_Y6_N29
\R.aluOp.ALUOpXor\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.aluOp.ALUOpXor_OTERM355\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluOp.ALUOpXor~q\);

-- Location: LABCELL_X73_Y6_N21
\R.aluOp.ALUOpXor_NEW354\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.aluOp.ALUOpXor_OTERM355\ = ( \vAluSrc2~0_combout\ & ( \Mux23~1_combout\ ) ) # ( !\vAluSrc2~0_combout\ & ( \R.aluOp.ALUOpXor~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111000000001111111100001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Mux23~1_combout\,
	datad => \ALT_INV_R.aluOp.ALUOpXor~q\,
	dataf => \ALT_INV_vAluSrc2~0_combout\,
	combout => \R.aluOp.ALUOpXor_OTERM355\);

-- Location: FF_X77_Y6_N2
\R.aluOp.ALUOpOr\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.aluOp.ALUOpOr_OTERM353\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluOp.ALUOpOr~q\);

-- Location: LABCELL_X77_Y6_N15
\Mux22~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux22~0_combout\ = ( \R.curInst\(13) & ( (!\Mux21~0_combout\ & (\R.curInst\(6) & ((\R.aluOp.ALUOpOr~q\)))) # (\Mux21~0_combout\ & ((!\R.curInst\(12)) # ((\R.curInst\(6) & \R.aluOp.ALUOpOr~q\)))) ) ) # ( !\R.curInst\(13) & ( (\R.curInst\(6) & 
-- \R.aluOp.ALUOpOr~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110011000000000011001101010000011100110101000001110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux21~0_combout\,
	datab => \ALT_INV_R.curInst\(6),
	datac => \ALT_INV_R.curInst\(12),
	datad => \ALT_INV_R.aluOp.ALUOpOr~q\,
	dataf => \ALT_INV_R.curInst\(13),
	combout => \Mux22~0_combout\);

-- Location: LABCELL_X77_Y6_N45
\Mux22~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux22~1_combout\ = ( \R.aluOp.ALUOpOr~q\ & ( \Mux22~0_combout\ & ( ((!\R.curInst\(3) & (!\Mux26~0_combout\)) # (\R.curInst\(3) & ((!\Mux123~0_combout\)))) # (\R.curInst\(4)) ) ) ) # ( !\R.aluOp.ALUOpOr~q\ & ( \Mux22~0_combout\ & ( (\R.curInst\(4) & 
-- !\R.curInst\(3)) ) ) ) # ( \R.aluOp.ALUOpOr~q\ & ( !\Mux22~0_combout\ & ( (!\R.curInst\(4) & ((!\R.curInst\(3) & (!\Mux26~0_combout\)) # (\R.curInst\(3) & ((!\Mux123~0_combout\))))) # (\R.curInst\(4) & (((\R.curInst\(3))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000100010001111010101010101000000001101110111110101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(4),
	datab => \ALT_INV_Mux26~0_combout\,
	datac => \ALT_INV_Mux123~0_combout\,
	datad => \ALT_INV_R.curInst\(3),
	datae => \ALT_INV_R.aluOp.ALUOpOr~q\,
	dataf => \ALT_INV_Mux22~0_combout\,
	combout => \Mux22~1_combout\);

-- Location: LABCELL_X77_Y6_N6
\R.aluOp.ALUOpOr_NEW352\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.aluOp.ALUOpOr_OTERM353\ = ( \vAluSrc2~0_combout\ & ( \Mux22~1_combout\ ) ) # ( !\vAluSrc2~0_combout\ & ( \R.aluOp.ALUOpOr~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100000000111111110000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluOp.ALUOpOr~q\,
	datad => \ALT_INV_Mux22~1_combout\,
	dataf => \ALT_INV_vAluSrc2~0_combout\,
	combout => \R.aluOp.ALUOpOr_OTERM353\);

-- Location: FF_X75_Y6_N47
\R.aluOp.ALUOpAnd\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.aluOp.ALUOpAnd_OTERM357\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluOp.ALUOpAnd~q\);

-- Location: FF_X75_Y6_N46
\R.aluOp.ALUOpAnd~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.aluOp.ALUOpAnd_OTERM357\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluOp.ALUOpAnd~DUPLICATE_q\);

-- Location: LABCELL_X77_Y6_N21
\Mux21~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux21~1_combout\ = ( \R.curInst\(13) & ( (!\Mux21~0_combout\ & (\R.curInst\(6) & (\R.aluOp.ALUOpAnd~q\))) # (\Mux21~0_combout\ & (((\R.curInst\(6) & \R.aluOp.ALUOpAnd~q\)) # (\R.curInst\(12)))) ) ) # ( !\R.curInst\(13) & ( (\R.curInst\(6) & 
-- \R.aluOp.ALUOpAnd~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000110000001100000011010101110000001101010111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux21~0_combout\,
	datab => \ALT_INV_R.curInst\(6),
	datac => \ALT_INV_R.aluOp.ALUOpAnd~q\,
	datad => \ALT_INV_R.curInst\(12),
	dataf => \ALT_INV_R.curInst\(13),
	combout => \Mux21~1_combout\);

-- Location: MLABCELL_X78_Y4_N0
\Mux21~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux21~2_combout\ = ( \Mux26~0_combout\ & ( \Mux21~1_combout\ & ( (!\R.curInst\(3) & (\R.curInst\(4))) # (\R.curInst\(3) & (\R.aluOp.ALUOpAnd~DUPLICATE_q\ & ((!\Mux123~0_combout\) # (\R.curInst\(4))))) ) ) ) # ( !\Mux26~0_combout\ & ( \Mux21~1_combout\ & 
-- ( (!\R.curInst\(4) & (\R.aluOp.ALUOpAnd~DUPLICATE_q\ & ((!\R.curInst\(3)) # (!\Mux123~0_combout\)))) # (\R.curInst\(4) & ((!\R.curInst\(3)) # ((\R.aluOp.ALUOpAnd~DUPLICATE_q\)))) ) ) ) # ( \Mux26~0_combout\ & ( !\Mux21~1_combout\ & ( (\R.curInst\(3) & 
-- (\R.aluOp.ALUOpAnd~DUPLICATE_q\ & ((!\Mux123~0_combout\) # (\R.curInst\(4))))) ) ) ) # ( !\Mux26~0_combout\ & ( !\Mux21~1_combout\ & ( (\R.aluOp.ALUOpAnd~DUPLICATE_q\ & ((!\R.curInst\(4) & ((!\R.curInst\(3)) # (!\Mux123~0_combout\))) # (\R.curInst\(4) & 
-- (\R.curInst\(3))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101100001001000000110000000101001111010011010100011101000101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(4),
	datab => \ALT_INV_R.curInst\(3),
	datac => \ALT_INV_R.aluOp.ALUOpAnd~DUPLICATE_q\,
	datad => \ALT_INV_Mux123~0_combout\,
	datae => \ALT_INV_Mux26~0_combout\,
	dataf => \ALT_INV_Mux21~1_combout\,
	combout => \Mux21~2_combout\);

-- Location: LABCELL_X75_Y6_N54
\R.aluOp.ALUOpAnd_NEW356\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.aluOp.ALUOpAnd_OTERM357\ = ( \Mux21~2_combout\ & ( (\R.aluOp.ALUOpAnd~q\) # (\vAluSrc2~0_combout\) ) ) # ( !\Mux21~2_combout\ & ( (!\vAluSrc2~0_combout\ & \R.aluOp.ALUOpAnd~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011110000000000001111000000001111111111110000111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_vAluSrc2~0_combout\,
	datad => \ALT_INV_R.aluOp.ALUOpAnd~q\,
	dataf => \ALT_INV_Mux21~2_combout\,
	combout => \R.aluOp.ALUOpAnd_OTERM357\);

-- Location: LABCELL_X71_Y7_N21
\Selector29~0_RTM0409\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector29~0_RTM0409_combout\ = ( \R.aluOp.ALUOpAnd_OTERM357\ & ( (!\Mux251~0_combout\ & (\NxR.aluData2[3]~18_combout\ & ((\R.aluOp.ALUOpOr_OTERM353\) # (\R.aluOp.ALUOpXor_OTERM355\)))) # (\Mux251~0_combout\ & (((\NxR.aluData2[3]~18_combout\) # 
-- (\R.aluOp.ALUOpOr_OTERM353\)) # (\R.aluOp.ALUOpXor_OTERM355\))) ) ) # ( !\R.aluOp.ALUOpAnd_OTERM357\ & ( (!\R.aluOp.ALUOpOr_OTERM353\ & (\R.aluOp.ALUOpXor_OTERM355\ & (!\Mux251~0_combout\ $ (!\NxR.aluData2[3]~18_combout\)))) # (\R.aluOp.ALUOpOr_OTERM353\ 
-- & (((\NxR.aluData2[3]~18_combout\) # (\Mux251~0_combout\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000011101110011000001110111001100000111011111110000011101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpXor_OTERM355\,
	datab => \ALT_INV_R.aluOp.ALUOpOr_OTERM353\,
	datac => \ALT_INV_Mux251~0_combout\,
	datad => \ALT_INV_NxR.aluData2[3]~18_combout\,
	dataf => \ALT_INV_R.aluOp.ALUOpAnd_OTERM357\,
	combout => \Selector29~0_RTM0409_combout\);

-- Location: FF_X71_Y7_N22
\Selector29~0_NEW_REG406\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector29~0_RTM0409_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector29~0_OTERM407\);

-- Location: LABCELL_X75_Y7_N0
\Selector29~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector29~1_combout\ = ( !\Selector29~0_OTERM407\ & ( \Selector32~3_OTERM379\ & ( !\ShiftLeft0~3_OTERM223\ ) ) ) # ( !\Selector29~0_OTERM407\ & ( !\Selector32~3_OTERM379\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111000000000000000011001100110011000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_ShiftLeft0~3_OTERM223\,
	datae => \ALT_INV_Selector29~0_OTERM407\,
	dataf => \ALT_INV_Selector32~3_OTERM379\,
	combout => \Selector29~1_combout\);

-- Location: LABCELL_X75_Y4_N0
\Mux149~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux149~0_combout\ = ( \R.curInst\(6) & ( (\R.curInst\(5) & (\R.curInst\(2) & (\R.curInst\(3) & !\R.curInst\(4)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000001000000000000000100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(5),
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_R.curInst\(3),
	datad => \ALT_INV_R.curInst\(4),
	dataf => \ALT_INV_R.curInst\(6),
	combout => \Mux149~0_combout\);

-- Location: LABCELL_X75_Y4_N36
\Mux123~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux123~2_combout\ = ( !\R.curInst\(4) & ( \R.curInst\(31) & ( (!\R.curInst\(3) & ((!\R.curInst\(6) & ((!\R.curInst\(2)))) # (\R.curInst\(6) & (\R.curInst\(5))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000010001010000000100000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(3),
	datab => \ALT_INV_R.curInst\(6),
	datac => \ALT_INV_R.curInst\(5),
	datad => \ALT_INV_R.curInst\(2),
	datae => \ALT_INV_R.curInst\(4),
	dataf => \ALT_INV_R.curInst\(31),
	combout => \Mux123~2_combout\);

-- Location: LABCELL_X75_Y4_N24
\Mux141~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux141~0_combout\ = ( \Mux123~2_combout\ & ( \R.curInst\(13) ) ) # ( !\Mux123~2_combout\ & ( \R.curInst\(13) & ( ((\vAluSrc1~0_combout\ & ((\R.curInst\(2)) # (\Mux124~0_combout\)))) # (\Mux149~0_combout\) ) ) ) # ( \Mux123~2_combout\ & ( !\R.curInst\(13) 
-- ) ) # ( !\Mux123~2_combout\ & ( !\R.curInst\(13) & ( (\Mux124~0_combout\ & \vAluSrc1~0_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010101111111111111111100001111011111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux124~0_combout\,
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_Mux149~0_combout\,
	datad => \ALT_INV_vAluSrc1~0_combout\,
	datae => \ALT_INV_Mux123~2_combout\,
	dataf => \ALT_INV_R.curInst\(13),
	combout => \Mux141~0_combout\);

-- Location: LABCELL_X77_Y1_N30
\Mux144~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux144~0_combout\ = ( \R.curInst\(5) & ( \R.curInst\(30) & ( (!\R.curInst\(4) & ((!\R.curInst\(2) & ((!\R.curInst\(3)))) # (\R.curInst\(2) & (\R.curInst\(6))))) ) ) ) # ( !\R.curInst\(5) & ( \R.curInst\(30) & ( (!\R.curInst\(6) & (!\R.curInst\(2) & 
-- !\R.curInst\(3))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000010100000000000001100010000000100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(6),
	datab => \ALT_INV_R.curInst\(4),
	datac => \ALT_INV_R.curInst\(2),
	datad => \ALT_INV_R.curInst\(3),
	datae => \ALT_INV_R.curInst\(5),
	dataf => \ALT_INV_R.curInst\(30),
	combout => \Mux144~0_combout\);

-- Location: LABCELL_X74_Y4_N9
\Mux130~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux130~0_combout\ = ( \Mux123~1_combout\ ) # ( !\Mux123~1_combout\ & ( (\vAluSrc1~0_combout\ & (((\R.curInst\(2) & \R.curInst\(24))) # (\Mux124~0_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000111000001010000011111111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux124~0_combout\,
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_vAluSrc1~0_combout\,
	datad => \ALT_INV_R.curInst\(24),
	dataf => \ALT_INV_Mux123~1_combout\,
	combout => \Mux130~0_combout\);

-- Location: FF_X74_Y7_N52
\Add2~33_OTERM719_NEW_REG824\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux246~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Add2~33_OTERM719_OTERM825\);

-- Location: LABCELL_X75_Y5_N36
\Mux146~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux146~0_combout\ = ( \R.curInst\(2) & ( \R.curInst\(5) & ( (!\R.curInst\(4) & (\R.curInst\(28) & \R.curInst\(6))) ) ) ) # ( !\R.curInst\(2) & ( \R.curInst\(5) & ( (!\R.curInst\(4) & (\R.curInst\(28) & !\R.curInst\(3))) ) ) ) # ( !\R.curInst\(2) & ( 
-- !\R.curInst\(5) & ( (\R.curInst\(28) & (!\R.curInst\(3) & !\R.curInst\(6))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011000000000000000000000000000000100000001000000000000000100010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(4),
	datab => \ALT_INV_R.curInst\(28),
	datac => \ALT_INV_R.curInst\(3),
	datad => \ALT_INV_R.curInst\(6),
	datae => \ALT_INV_R.curInst\(2),
	dataf => \ALT_INV_R.curInst\(5),
	combout => \Mux146~0_combout\);

-- Location: LABCELL_X77_Y1_N9
\Mux147~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux147~0_combout\ = ( \R.curInst\(27) & ( \R.curInst\(5) & ( (!\R.curInst\(4) & ((!\R.curInst\(2) & (!\R.curInst\(3))) # (\R.curInst\(2) & ((\R.curInst\(6)))))) ) ) ) # ( \R.curInst\(27) & ( !\R.curInst\(5) & ( (!\R.curInst\(2) & (!\R.curInst\(3) & 
-- !\R.curInst\(6))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000100010000000000000000000000000001000000011010000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(2),
	datab => \ALT_INV_R.curInst\(3),
	datac => \ALT_INV_R.curInst\(4),
	datad => \ALT_INV_R.curInst\(6),
	datae => \ALT_INV_R.curInst\(27),
	dataf => \ALT_INV_R.curInst\(5),
	combout => \Mux147~0_combout\);

-- Location: FF_X73_Y5_N2
\R.aluData1[29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Mux225~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData1\(29));

-- Location: MLABCELL_X72_Y5_N18
\Selector17~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector17~0_combout\ = ( \R.aluOp.ALUOpSRA_OTERM363\ & ( (\NxR.aluData2[4]~20_combout\ & \Mux223~0_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000011110000000000001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_NxR.aluData2[4]~20_combout\,
	datad => \ALT_INV_Mux223~0_combout\,
	dataf => \ALT_INV_R.aluOp.ALUOpSRA_OTERM363\,
	combout => \Selector17~0_combout\);

-- Location: FF_X72_Y5_N19
\Selector17~0_NEW_REG390\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector17~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector17~0_OTERM391\);

-- Location: LABCELL_X74_Y4_N6
\Mux125~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux125~0_combout\ = ( \Mux123~1_combout\ ) # ( !\Mux123~1_combout\ & ( (\vAluSrc1~0_combout\ & (((\R.curInst\(2) & \R.curInst\(29))) # (\Mux124~0_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010111000000000101011111111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux124~0_combout\,
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_R.curInst\(29),
	datad => \ALT_INV_vAluSrc1~0_combout\,
	dataf => \ALT_INV_Mux123~1_combout\,
	combout => \Mux125~0_combout\);

-- Location: LABCELL_X81_Y5_N48
\Add0~105\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~105_sumout\ = SUM(( \R.curPC\(28) ) + ( GND ) + ( \Add0~102\ ))
-- \Add0~106\ = CARRY(( \R.curPC\(28) ) + ( GND ) + ( \Add0~102\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.curPC\(28),
	cin => \Add0~102\,
	sumout => \Add0~105_sumout\,
	cout => \Add0~106\);

-- Location: LABCELL_X81_Y5_N51
\Add0~109\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~109_sumout\ = SUM(( \R.curPC\(29) ) + ( GND ) + ( \Add0~106\ ))
-- \Add0~110\ = CARRY(( \R.curPC\(29) ) + ( GND ) + ( \Add0~106\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curPC\(29),
	cin => \Add0~106\,
	sumout => \Add0~109_sumout\,
	cout => \Add0~110\);

-- Location: FF_X67_Y8_N56
\RegFile[13][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(27),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][27]~q\);

-- Location: MLABCELL_X72_Y8_N9
\RegFile[15][27]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[15][27]~feeder_combout\ = ( \R.regWriteData\(27) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(27),
	combout => \RegFile[15][27]~feeder_combout\);

-- Location: FF_X72_Y8_N10
\RegFile[15][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[15][27]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][27]~q\);

-- Location: LABCELL_X67_Y8_N33
\RegFile[14][27]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[14][27]~feeder_combout\ = ( \R.regWriteData\(27) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(27),
	combout => \RegFile[14][27]~feeder_combout\);

-- Location: FF_X67_Y8_N35
\RegFile[14][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[14][27]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][27]~q\);

-- Location: FF_X67_Y8_N2
\RegFile[9][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(27),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][27]~q\);

-- Location: FF_X64_Y8_N1
\RegFile[11][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(27),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][27]~q\);

-- Location: FF_X64_Y8_N19
\RegFile[10][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(27),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][27]~q\);

-- Location: FF_X66_Y5_N46
\RegFile[8][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(27),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][27]~q\);

-- Location: LABCELL_X67_Y8_N39
\Mux63~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux63~14_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[8][27]~q\))) # (\R.curInst\(15) & (\RegFile[9][27]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[10][27]~q\))) # (\R.curInst\(15) & (\RegFile[11][27]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][27]~q\,
	datab => \ALT_INV_RegFile[11][27]~q\,
	datac => \ALT_INV_RegFile[10][27]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][27]~q\,
	combout => \Mux63~14_combout\);

-- Location: FF_X74_Y8_N28
\RegFile[12][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(27),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][27]~q\);

-- Location: LABCELL_X67_Y8_N54
\Mux63~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux63~1_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux63~14_combout\)))) # (\R.curInst\(17) & ((!\Mux63~14_combout\ & ((\RegFile[12][27]~q\))) # (\Mux63~14_combout\ & (\RegFile[13][27]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux63~14_combout\)))) # (\R.curInst\(17) & ((!\Mux63~14_combout\ & ((\RegFile[14][27]~q\))) # (\Mux63~14_combout\ & (\RegFile[15][27]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][27]~q\,
	datab => \ALT_INV_RegFile[15][27]~q\,
	datac => \ALT_INV_RegFile[14][27]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux63~14_combout\,
	datag => \ALT_INV_RegFile[12][27]~q\,
	combout => \Mux63~1_combout\);

-- Location: FF_X70_Y7_N8
\RegFile[23][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(27),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][27]~q\);

-- Location: LABCELL_X73_Y10_N51
\RegFile[22][27]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[22][27]~feeder_combout\ = ( \R.regWriteData\(27) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(27),
	combout => \RegFile[22][27]~feeder_combout\);

-- Location: FF_X73_Y10_N52
\RegFile[22][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[22][27]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][27]~q\);

-- Location: LABCELL_X70_Y7_N54
\RegFile[21][27]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[21][27]~feeder_combout\ = ( \R.regWriteData\(27) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(27),
	combout => \RegFile[21][27]~feeder_combout\);

-- Location: FF_X70_Y7_N55
\RegFile[21][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[21][27]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][27]~q\);

-- Location: FF_X66_Y4_N8
\RegFile[17][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(27),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][27]~q\);

-- Location: LABCELL_X66_Y4_N39
\RegFile[18][27]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[18][27]~feeder_combout\ = ( \R.regWriteData\(27) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(27),
	combout => \RegFile[18][27]~feeder_combout\);

-- Location: FF_X66_Y4_N41
\RegFile[18][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][27]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][27]~q\);

-- Location: LABCELL_X66_Y4_N57
\RegFile[19][27]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[19][27]~feeder_combout\ = ( \R.regWriteData\(27) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(27),
	combout => \RegFile[19][27]~feeder_combout\);

-- Location: FF_X66_Y4_N58
\RegFile[19][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[19][27]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][27]~q\);

-- Location: LABCELL_X61_Y8_N6
\RegFile[16][27]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[16][27]~feeder_combout\ = ( \R.regWriteData\(27) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(27),
	combout => \RegFile[16][27]~feeder_combout\);

-- Location: FF_X61_Y8_N7
\RegFile[16][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[16][27]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][27]~q\);

-- Location: LABCELL_X70_Y4_N48
\Mux63~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux63~18_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[16][27]~q\))) # (\R.curInst\(15) & (\RegFile[17][27]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & (\RegFile[18][27]~q\)) # (\R.curInst\(15) & ((\RegFile[19][27]~q\)))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001110111011101110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[17][27]~q\,
	datac => \ALT_INV_RegFile[18][27]~q\,
	datad => \ALT_INV_RegFile[19][27]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][27]~q\,
	combout => \Mux63~18_combout\);

-- Location: FF_X68_Y6_N8
\RegFile[20][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(27),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][27]~q\);

-- Location: LABCELL_X70_Y7_N6
\Mux63~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux63~5_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux63~18_combout\))))) # (\R.curInst\(17) & (((!\Mux63~18_combout\ & (\RegFile[20][27]~q\)) # (\Mux63~18_combout\ & ((\RegFile[21][27]~q\)))))) ) ) # ( \R.curInst\(16) & ( 
-- (!\R.curInst\(17) & ((((\Mux63~18_combout\))))) # (\R.curInst\(17) & (((!\Mux63~18_combout\ & ((\RegFile[22][27]~q\))) # (\Mux63~18_combout\ & (\RegFile[23][27]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110101010111111111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[23][27]~q\,
	datac => \ALT_INV_RegFile[22][27]~q\,
	datad => \ALT_INV_RegFile[21][27]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux63~18_combout\,
	datag => \ALT_INV_RegFile[20][27]~q\,
	combout => \Mux63~5_combout\);

-- Location: FF_X67_Y5_N13
\RegFile[4][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(27),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][27]~q\);

-- Location: FF_X65_Y6_N20
\RegFile[6][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(27),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][27]~q\);

-- Location: MLABCELL_X59_Y6_N3
\RegFile[5][27]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[5][27]~feeder_combout\ = ( \R.regWriteData\(27) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(27),
	combout => \RegFile[5][27]~feeder_combout\);

-- Location: FF_X59_Y6_N4
\RegFile[5][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[5][27]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][27]~q\);

-- Location: FF_X65_Y6_N50
\RegFile[7][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(27),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][27]~q\);

-- Location: MLABCELL_X65_Y6_N48
\Mux63~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux63~0_combout\ = ( \RegFile[7][27]~q\ & ( \R.curInst\(15) & ( (\RegFile[5][27]~q\) # (\R.curInst\(16)) ) ) ) # ( !\RegFile[7][27]~q\ & ( \R.curInst\(15) & ( (!\R.curInst\(16) & \RegFile[5][27]~q\) ) ) ) # ( \RegFile[7][27]~q\ & ( !\R.curInst\(15) & ( 
-- (!\R.curInst\(16) & (\RegFile[4][27]~q\)) # (\R.curInst\(16) & ((\RegFile[6][27]~q\))) ) ) ) # ( !\RegFile[7][27]~q\ & ( !\R.curInst\(15) & ( (!\R.curInst\(16) & (\RegFile[4][27]~q\)) # (\R.curInst\(16) & ((\RegFile[6][27]~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100011101000111010001110100011100000000110011000011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[4][27]~q\,
	datab => \ALT_INV_R.curInst\(16),
	datac => \ALT_INV_RegFile[6][27]~q\,
	datad => \ALT_INV_RegFile[5][27]~q\,
	datae => \ALT_INV_RegFile[7][27]~q\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux63~0_combout\);

-- Location: LABCELL_X70_Y7_N48
\RegFile[3][27]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[3][27]~feeder_combout\ = ( \R.regWriteData\(27) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(27),
	combout => \RegFile[3][27]~feeder_combout\);

-- Location: FF_X70_Y7_N50
\RegFile[3][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[3][27]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][27]~q\);

-- Location: FF_X65_Y6_N14
\RegFile[2][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(27),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][27]~q\);

-- Location: MLABCELL_X59_Y6_N42
\RegFile[1][27]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[1][27]~feeder_combout\ = ( \R.regWriteData\(27) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(27),
	combout => \RegFile[1][27]~feeder_combout\);

-- Location: FF_X59_Y6_N43
\RegFile[1][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[1][27]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][27]~q\);

-- Location: MLABCELL_X65_Y6_N12
\Mux63~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux63~26_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\RegFile[1][27]~q\ & \R.curInst\(15))))) # (\R.curInst\(17) & (\Mux63~0_combout\))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[2][27]~q\))) # 
-- (\R.curInst\(15) & (\RegFile[3][27]~q\))))) # (\R.curInst\(17) & (\Mux63~0_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000001010101000011110101010100001111010101010011001101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux63~0_combout\,
	datab => \ALT_INV_RegFile[3][27]~q\,
	datac => \ALT_INV_RegFile[2][27]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[1][27]~q\,
	combout => \Mux63~26_combout\);

-- Location: FF_X73_Y5_N50
\RegFile[31][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(27),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][27]~q\);

-- Location: LABCELL_X70_Y9_N12
\RegFile[30][27]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[30][27]~feeder_combout\ = ( \R.regWriteData\(27) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(27),
	combout => \RegFile[30][27]~feeder_combout\);

-- Location: FF_X70_Y9_N13
\RegFile[30][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[30][27]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][27]~q\);

-- Location: FF_X67_Y4_N38
\RegFile[27][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(27),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][27]~q\);

-- Location: FF_X71_Y4_N50
\RegFile[25][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(27),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][27]~q\);

-- Location: LABCELL_X67_Y4_N54
\RegFile[26][27]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[26][27]~feeder_combout\ = \R.regWriteData\(27)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.regWriteData\(27),
	combout => \RegFile[26][27]~feeder_combout\);

-- Location: FF_X67_Y4_N56
\RegFile[26][27]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[26][27]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][27]~DUPLICATE_q\);

-- Location: LABCELL_X56_Y4_N0
\RegFile[24][27]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[24][27]~feeder_combout\ = ( \R.regWriteData\(27) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(27),
	combout => \RegFile[24][27]~feeder_combout\);

-- Location: FF_X56_Y4_N1
\RegFile[24][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[24][27]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][27]~q\);

-- Location: LABCELL_X67_Y4_N36
\Mux63~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux63~22_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[24][27]~q\))) # (\R.curInst\(15) & (\RegFile[25][27]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[26][27]~DUPLICATE_q\))) # (\R.curInst\(15) & (\RegFile[27][27]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[27][27]~q\,
	datab => \ALT_INV_RegFile[25][27]~q\,
	datac => \ALT_INV_RegFile[26][27]~DUPLICATE_q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][27]~q\,
	combout => \Mux63~22_combout\);

-- Location: FF_X74_Y8_N58
\RegFile[28][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(27),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][27]~q\);

-- Location: LABCELL_X73_Y5_N48
\Mux63~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux63~9_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux63~22_combout\)))) # (\R.curInst\(17) & ((!\Mux63~22_combout\ & ((\RegFile[28][27]~q\))) # (\Mux63~22_combout\ & (\RegFile[29][27]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux63~22_combout\)))) # (\R.curInst\(17) & ((!\Mux63~22_combout\ & ((\RegFile[30][27]~q\))) # (\Mux63~22_combout\ & (\RegFile[31][27]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][27]~q\,
	datab => \ALT_INV_RegFile[29][27]~q\,
	datac => \ALT_INV_RegFile[30][27]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux63~22_combout\,
	datag => \ALT_INV_RegFile[28][27]~q\,
	combout => \Mux63~9_combout\);

-- Location: LABCELL_X73_Y4_N48
\Mux63~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux63~13_combout\ = ( \Mux63~26_combout\ & ( \Mux63~9_combout\ & ( (!\R.curInst\(19) & ((!\R.curInst\(18)) # ((\Mux63~1_combout\)))) # (\R.curInst\(19) & (((\Mux63~5_combout\)) # (\R.curInst\(18)))) ) ) ) # ( !\Mux63~26_combout\ & ( \Mux63~9_combout\ & ( 
-- (!\R.curInst\(19) & (\R.curInst\(18) & (\Mux63~1_combout\))) # (\R.curInst\(19) & (((\Mux63~5_combout\)) # (\R.curInst\(18)))) ) ) ) # ( \Mux63~26_combout\ & ( !\Mux63~9_combout\ & ( (!\R.curInst\(19) & ((!\R.curInst\(18)) # ((\Mux63~1_combout\)))) # 
-- (\R.curInst\(19) & (!\R.curInst\(18) & ((\Mux63~5_combout\)))) ) ) ) # ( !\Mux63~26_combout\ & ( !\Mux63~9_combout\ & ( (!\R.curInst\(19) & (\R.curInst\(18) & (\Mux63~1_combout\))) # (\R.curInst\(19) & (!\R.curInst\(18) & ((\Mux63~5_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001001000110100010101100111000010011010101111001101111011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(19),
	datab => \ALT_INV_R.curInst\(18),
	datac => \ALT_INV_Mux63~1_combout\,
	datad => \ALT_INV_Mux63~5_combout\,
	datae => \ALT_INV_Mux63~26_combout\,
	dataf => \ALT_INV_Mux63~9_combout\,
	combout => \Mux63~13_combout\);

-- Location: LABCELL_X73_Y4_N45
\Mux227~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux227~0_combout\ = ( \Mux63~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC\(27)))) ) ) # ( !\Mux63~13_combout\ & ( (\vAluSrc1~2_combout\ & (!\vAluSrc1~1_combout\ & \R.curPC\(27))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001000100000000000100010010001000110011001000100011001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluSrc1~2_combout\,
	datab => \ALT_INV_vAluSrc1~1_combout\,
	datad => \ALT_INV_R.curPC\(27),
	dataf => \ALT_INV_Mux63~13_combout\,
	combout => \Mux227~0_combout\);

-- Location: FF_X73_Y4_N40
\R.aluData1[27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux227~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData1\(27));

-- Location: LABCELL_X75_Y4_N18
\Mux128~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux128~0_combout\ = ( \vAluSrc1~0_combout\ & ( (((\R.curInst\(2) & \R.curInst\(26))) # (\Mux123~1_combout\)) # (\Mux124~0_combout\) ) ) # ( !\vAluSrc1~0_combout\ & ( \Mux123~1_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111000000001111111101010111111111110101011111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux124~0_combout\,
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_R.curInst\(26),
	datad => \ALT_INV_Mux123~1_combout\,
	dataf => \ALT_INV_vAluSrc1~0_combout\,
	combout => \Mux128~0_combout\);

-- Location: FF_X67_Y7_N14
\RegFile[3][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(26),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][26]~q\);

-- Location: FF_X60_Y4_N41
\RegFile[2][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(26),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][26]~q\);

-- Location: FF_X61_Y4_N49
\RegFile[7][26]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(26),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][26]~DUPLICATE_q\);

-- Location: FF_X61_Y4_N8
\RegFile[6][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(26),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][26]~q\);

-- Location: LABCELL_X62_Y8_N48
\RegFile[5][26]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[5][26]~feeder_combout\ = ( \R.regWriteData\(26) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(26),
	combout => \RegFile[5][26]~feeder_combout\);

-- Location: FF_X62_Y8_N49
\RegFile[5][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[5][26]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][26]~q\);

-- Location: LABCELL_X56_Y4_N39
\RegFile[4][26]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[4][26]~feeder_combout\ = ( \R.regWriteData\(26) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(26),
	combout => \RegFile[4][26]~feeder_combout\);

-- Location: FF_X56_Y4_N40
\RegFile[4][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[4][26]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][26]~q\);

-- Location: LABCELL_X67_Y4_N15
\Mux96~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux96~0_combout\ = ( \R.curInst\(21) & ( \R.curInst\(20) & ( \RegFile[7][26]~DUPLICATE_q\ ) ) ) # ( !\R.curInst\(21) & ( \R.curInst\(20) & ( \RegFile[5][26]~q\ ) ) ) # ( \R.curInst\(21) & ( !\R.curInst\(20) & ( \RegFile[6][26]~q\ ) ) ) # ( 
-- !\R.curInst\(21) & ( !\R.curInst\(20) & ( \RegFile[4][26]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111001100110011001100001111000011110101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[7][26]~DUPLICATE_q\,
	datab => \ALT_INV_RegFile[6][26]~q\,
	datac => \ALT_INV_RegFile[5][26]~q\,
	datad => \ALT_INV_RegFile[4][26]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	combout => \Mux96~0_combout\);

-- Location: LABCELL_X61_Y5_N15
\RegFile[1][26]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[1][26]~feeder_combout\ = ( \R.regWriteData\(26) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(26),
	combout => \RegFile[1][26]~feeder_combout\);

-- Location: FF_X61_Y5_N16
\RegFile[1][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[1][26]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][26]~q\);

-- Location: LABCELL_X67_Y7_N12
\Mux96~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux96~26_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (\R.curInst\(20) & (\RegFile[1][26]~q\))) # (\R.curInst\(22) & (((\Mux96~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (((\RegFile[2][26]~q\)))) # 
-- (\R.curInst\(20) & (\RegFile[3][26]~q\)))) # (\R.curInst\(22) & ((((\Mux96~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000000000110110000000000000101111111110001101111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(20),
	datab => \ALT_INV_RegFile[3][26]~q\,
	datac => \ALT_INV_RegFile[2][26]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux96~0_combout\,
	datag => \ALT_INV_RegFile[1][26]~q\,
	combout => \Mux96~26_combout\);

-- Location: FF_X73_Y4_N26
\RegFile[23][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(26),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][26]~q\);

-- Location: FF_X72_Y9_N52
\RegFile[22][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(26),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][26]~q\);

-- Location: FF_X70_Y4_N32
\RegFile[17][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(26),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][26]~q\);

-- Location: LABCELL_X71_Y4_N42
\RegFile[18][26]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[18][26]~feeder_combout\ = ( \R.regWriteData\(26) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(26),
	combout => \RegFile[18][26]~feeder_combout\);

-- Location: FF_X71_Y4_N43
\RegFile[18][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][26]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][26]~q\);

-- Location: FF_X70_Y4_N8
\RegFile[19][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(26),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][26]~q\);

-- Location: LABCELL_X63_Y9_N57
\RegFile[16][26]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[16][26]~feeder_combout\ = ( \R.regWriteData\(26) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(26),
	combout => \RegFile[16][26]~feeder_combout\);

-- Location: FF_X63_Y9_N58
\RegFile[16][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[16][26]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][26]~q\);

-- Location: LABCELL_X70_Y4_N30
\Mux96~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux96~18_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[16][26]~q\))) # (\R.curInst\(20) & (\RegFile[17][26]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & (\RegFile[18][26]~q\)) # (\R.curInst\(20) & ((\RegFile[19][26]~q\)))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001110111011101110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[17][26]~q\,
	datac => \ALT_INV_RegFile[18][26]~q\,
	datad => \ALT_INV_RegFile[19][26]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][26]~q\,
	combout => \Mux96~18_combout\);

-- Location: FF_X77_Y8_N40
\RegFile[20][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(26),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][26]~q\);

-- Location: LABCELL_X70_Y6_N42
\Mux96~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux96~5_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux96~18_combout\)))) # (\R.curInst\(22) & ((!\Mux96~18_combout\ & ((\RegFile[20][26]~q\))) # (\Mux96~18_combout\ & (\RegFile[21][26]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux96~18_combout\)))) # (\R.curInst\(22) & ((!\Mux96~18_combout\ & ((\RegFile[22][26]~q\))) # (\Mux96~18_combout\ & (\RegFile[23][26]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][26]~q\,
	datab => \ALT_INV_RegFile[23][26]~q\,
	datac => \ALT_INV_RegFile[22][26]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux96~18_combout\,
	datag => \ALT_INV_RegFile[20][26]~q\,
	combout => \Mux96~5_combout\);

-- Location: FF_X71_Y4_N2
\RegFile[29][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(26),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][26]~q\);

-- Location: LABCELL_X73_Y8_N54
\RegFile[30][26]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[30][26]~feeder_combout\ = ( \R.regWriteData\(26) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(26),
	combout => \RegFile[30][26]~feeder_combout\);

-- Location: FF_X73_Y8_N55
\RegFile[30][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[30][26]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][26]~q\);

-- Location: FF_X73_Y4_N56
\RegFile[31][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(26),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][26]~q\);

-- Location: FF_X71_Y4_N35
\RegFile[25][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(26),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][26]~q\);

-- Location: LABCELL_X67_Y4_N57
\RegFile[26][26]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[26][26]~feeder_combout\ = ( \R.regWriteData\(26) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(26),
	combout => \RegFile[26][26]~feeder_combout\);

-- Location: FF_X67_Y4_N58
\RegFile[26][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[26][26]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][26]~q\);

-- Location: FF_X67_Y4_N44
\RegFile[27][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(26),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][26]~q\);

-- Location: LABCELL_X57_Y4_N51
\RegFile[24][26]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[24][26]~feeder_combout\ = ( \R.regWriteData\(26) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(26),
	combout => \RegFile[24][26]~feeder_combout\);

-- Location: FF_X57_Y4_N52
\RegFile[24][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[24][26]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][26]~q\);

-- Location: LABCELL_X71_Y4_N33
\Mux96~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux96~22_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[24][26]~q\))) # (\R.curInst\(20) & (\RegFile[25][26]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & (\RegFile[26][26]~q\)) # (\R.curInst\(20) & ((\RegFile[27][26]~q\)))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001110111011101110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[25][26]~q\,
	datac => \ALT_INV_RegFile[26][26]~q\,
	datad => \ALT_INV_RegFile[27][26]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][26]~q\,
	combout => \Mux96~22_combout\);

-- Location: FF_X70_Y9_N1
\RegFile[28][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(26),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][26]~q\);

-- Location: LABCELL_X71_Y4_N0
\Mux96~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux96~9_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux96~22_combout\))))) # (\R.curInst\(22) & (((!\Mux96~22_combout\ & ((\RegFile[28][26]~q\))) # (\Mux96~22_combout\ & (\RegFile[29][26]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux96~22_combout\)))) # (\R.curInst\(22) & ((!\Mux96~22_combout\ & (\RegFile[30][26]~q\)) # (\Mux96~22_combout\ & ((\RegFile[31][26]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[29][26]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[30][26]~q\,
	datad => \ALT_INV_RegFile[31][26]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux96~22_combout\,
	datag => \ALT_INV_RegFile[28][26]~q\,
	combout => \Mux96~9_combout\);

-- Location: FF_X70_Y6_N14
\RegFile[15][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(26),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][26]~q\);

-- Location: LABCELL_X56_Y8_N9
\RegFile[14][26]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[14][26]~feeder_combout\ = ( \R.regWriteData\(26) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(26),
	combout => \RegFile[14][26]~feeder_combout\);

-- Location: FF_X56_Y8_N10
\RegFile[14][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[14][26]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][26]~q\);

-- Location: FF_X63_Y8_N20
\RegFile[13][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(26),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][26]~q\);

-- Location: FF_X64_Y8_N38
\RegFile[11][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(26),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][26]~q\);

-- Location: FF_X63_Y8_N8
\RegFile[9][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(26),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][26]~q\);

-- Location: FF_X64_Y8_N31
\RegFile[10][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(26),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][26]~q\);

-- Location: FF_X63_Y8_N34
\RegFile[8][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(26),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][26]~q\);

-- Location: LABCELL_X64_Y8_N36
\Mux96~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux96~14_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[8][26]~q\))) # (\R.curInst\(20) & (\RegFile[9][26]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[10][26]~q\))) # (\R.curInst\(20) & (\RegFile[11][26]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[11][26]~q\,
	datab => \ALT_INV_RegFile[9][26]~q\,
	datac => \ALT_INV_RegFile[10][26]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][26]~q\,
	combout => \Mux96~14_combout\);

-- Location: LABCELL_X66_Y10_N54
\RegFile[12][26]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[12][26]~feeder_combout\ = ( \R.regWriteData\(26) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(26),
	combout => \RegFile[12][26]~feeder_combout\);

-- Location: FF_X66_Y10_N55
\RegFile[12][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[12][26]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][26]~q\);

-- Location: LABCELL_X70_Y6_N12
\Mux96~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux96~1_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux96~14_combout\)))) # (\R.curInst\(22) & ((!\Mux96~14_combout\ & (\RegFile[12][26]~q\)) # (\Mux96~14_combout\ & ((\RegFile[13][26]~q\)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) 
-- & ((((\Mux96~14_combout\))))) # (\R.curInst\(22) & (((!\Mux96~14_combout\ & ((\RegFile[14][26]~q\))) # (\Mux96~14_combout\ & (\RegFile[15][26]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111001100111111111101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][26]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[14][26]~q\,
	datad => \ALT_INV_RegFile[13][26]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux96~14_combout\,
	datag => \ALT_INV_RegFile[12][26]~q\,
	combout => \Mux96~1_combout\);

-- Location: LABCELL_X70_Y6_N48
\Mux96~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux96~13_combout\ = ( \Mux96~9_combout\ & ( \Mux96~1_combout\ & ( ((!\R.curInst\(24) & (\Mux96~26_combout\)) # (\R.curInst\(24) & ((\Mux96~5_combout\)))) # (\R.curInst\(23)) ) ) ) # ( !\Mux96~9_combout\ & ( \Mux96~1_combout\ & ( (!\R.curInst\(24) & 
-- (((\Mux96~26_combout\)) # (\R.curInst\(23)))) # (\R.curInst\(24) & (!\R.curInst\(23) & ((\Mux96~5_combout\)))) ) ) ) # ( \Mux96~9_combout\ & ( !\Mux96~1_combout\ & ( (!\R.curInst\(24) & (!\R.curInst\(23) & (\Mux96~26_combout\))) # (\R.curInst\(24) & 
-- (((\Mux96~5_combout\)) # (\R.curInst\(23)))) ) ) ) # ( !\Mux96~9_combout\ & ( !\Mux96~1_combout\ & ( (!\R.curInst\(23) & ((!\R.curInst\(24) & (\Mux96~26_combout\)) # (\R.curInst\(24) & ((\Mux96~5_combout\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000100001001100000110010101110100101010011011100011101101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(24),
	datab => \ALT_INV_R.curInst\(23),
	datac => \ALT_INV_Mux96~26_combout\,
	datad => \ALT_INV_Mux96~5_combout\,
	datae => \ALT_INV_Mux96~9_combout\,
	dataf => \ALT_INV_Mux96~1_combout\,
	combout => \Mux96~13_combout\);

-- Location: LABCELL_X73_Y4_N3
\NxR.aluData2[26]~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[26]~25_combout\ = ( \Mux96~13_combout\ & ( (!\vAluSrc2~1_combout\) # ((\Equal4~1_combout\ & \Mux128~0_combout\)) ) ) # ( !\Mux96~13_combout\ & ( (\vAluSrc2~1_combout\ & (\Equal4~1_combout\ & \Mux128~0_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000010001000000000001000110101010101110111010101010111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluSrc2~1_combout\,
	datab => \ALT_INV_Equal4~1_combout\,
	datad => \ALT_INV_Mux128~0_combout\,
	dataf => \ALT_INV_Mux96~13_combout\,
	combout => \NxR.aluData2[26]~25_combout\);

-- Location: FF_X73_Y4_N35
\R.aluData2[26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \NxR.aluData2[26]~25_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData2\(26));

-- Location: FF_X73_Y4_N16
\R.aluData1[26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux228~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData1\(26));

-- Location: LABCELL_X81_Y5_N36
\Add0~89\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~89_sumout\ = SUM(( \R.curPC\(24) ) + ( GND ) + ( \Add0~86\ ))
-- \Add0~90\ = CARRY(( \R.curPC\(24) ) + ( GND ) + ( \Add0~86\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.curPC\(24),
	cin => \Add0~86\,
	sumout => \Add0~89_sumout\,
	cout => \Add0~90\);

-- Location: LABCELL_X81_Y5_N39
\Add0~93\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~93_sumout\ = SUM(( \R.curPC\(25) ) + ( GND ) + ( \Add0~90\ ))
-- \Add0~94\ = CARRY(( \R.curPC\(25) ) + ( GND ) + ( \Add0~90\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.curPC\(25),
	cin => \Add0~90\,
	sumout => \Add0~93_sumout\,
	cout => \Add0~94\);

-- Location: FF_X72_Y5_N29
\R.aluData1[31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux223~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData1\(31));

-- Location: LABCELL_X77_Y9_N54
\ShiftRight1~55\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~55_combout\ = ( \ShiftRight1~13_OTERM15\ & ( \R.aluData1\(31) & ( ((\R.aluData2\(2)) # (\R.aluData2\(3))) # (\ShiftRight1~12_OTERM57\) ) ) ) # ( !\ShiftRight1~13_OTERM15\ & ( \R.aluData1\(31) & ( ((\ShiftRight1~12_OTERM57\ & 
-- !\R.aluData2\(2))) # (\R.aluData2\(3)) ) ) ) # ( \ShiftRight1~13_OTERM15\ & ( !\R.aluData1\(31) & ( (!\R.aluData2\(3) & ((\R.aluData2\(2)) # (\ShiftRight1~12_OTERM57\))) ) ) ) # ( !\ShiftRight1~13_OTERM15\ & ( !\R.aluData1\(31) & ( 
-- (\ShiftRight1~12_OTERM57\ & (!\R.aluData2\(3) & !\R.aluData2\(2))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101000000000000010100001111000001011111000011110101111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~12_OTERM57\,
	datac => \ALT_INV_R.aluData2\(3),
	datad => \ALT_INV_R.aluData2\(2),
	datae => \ALT_INV_ShiftRight1~13_OTERM15\,
	dataf => \ALT_INV_R.aluData1\(31),
	combout => \ShiftRight1~55_combout\);

-- Location: LABCELL_X81_Y5_N54
\Add0~113\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~113_sumout\ = SUM(( \R.curPC[30]~DUPLICATE_q\ ) + ( GND ) + ( \Add0~110\ ))
-- \Add0~114\ = CARRY(( \R.curPC[30]~DUPLICATE_q\ ) + ( GND ) + ( \Add0~110\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.curPC[30]~DUPLICATE_q\,
	cin => \Add0~110\,
	sumout => \Add0~113_sumout\,
	cout => \Add0~114\);

-- Location: LABCELL_X74_Y4_N3
\Mux124~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux124~1_combout\ = ( \Mux124~0_combout\ & ( (\Mux123~1_combout\) # (\vAluSrc1~0_combout\) ) ) # ( !\Mux124~0_combout\ & ( ((\vAluSrc1~0_combout\ & (\R.curInst\(2) & \R.curInst\(30)))) # (\Mux123~1_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000111111111000000011111111101010101111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluSrc1~0_combout\,
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_R.curInst\(30),
	datad => \ALT_INV_Mux123~1_combout\,
	dataf => \ALT_INV_Mux124~0_combout\,
	combout => \Mux124~1_combout\);

-- Location: FF_X59_Y2_N22
\RegFile[29][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(30),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][30]~q\);

-- Location: LABCELL_X66_Y3_N54
\RegFile[30][30]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[30][30]~feeder_combout\ = ( \R.regWriteData\(30) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(30),
	combout => \RegFile[30][30]~feeder_combout\);

-- Location: FF_X66_Y3_N55
\RegFile[30][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[30][30]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][30]~q\);

-- Location: FF_X66_Y3_N32
\RegFile[31][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(30),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][30]~q\);

-- Location: LABCELL_X63_Y2_N42
\RegFile[27][30]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[27][30]~feeder_combout\ = ( \R.regWriteData\(30) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(30),
	combout => \RegFile[27][30]~feeder_combout\);

-- Location: FF_X63_Y2_N43
\RegFile[27][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[27][30]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][30]~q\);

-- Location: LABCELL_X60_Y2_N9
\RegFile[26][30]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[26][30]~feeder_combout\ = ( \R.regWriteData\(30) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(30),
	combout => \RegFile[26][30]~feeder_combout\);

-- Location: FF_X60_Y2_N10
\RegFile[26][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[26][30]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][30]~q\);

-- Location: FF_X63_Y2_N2
\RegFile[25][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(30),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][30]~q\);

-- Location: FF_X59_Y2_N53
\RegFile[24][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(30),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][30]~q\);

-- Location: LABCELL_X63_Y2_N0
\Mux92~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux92~22_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & (\RegFile[24][30]~q\)) # (\R.curInst\(20) & ((\RegFile[25][30]~q\)))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & ((\RegFile[26][30]~q\))) # (\R.curInst\(20) & (\RegFile[27][30]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001010101111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[27][30]~q\,
	datac => \ALT_INV_RegFile[26][30]~q\,
	datad => \ALT_INV_RegFile[25][30]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][30]~q\,
	combout => \Mux92~22_combout\);

-- Location: LABCELL_X66_Y3_N0
\RegFile[28][30]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[28][30]~feeder_combout\ = \R.regWriteData\(30)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.regWriteData\(30),
	combout => \RegFile[28][30]~feeder_combout\);

-- Location: FF_X66_Y3_N2
\RegFile[28][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[28][30]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][30]~q\);

-- Location: LABCELL_X62_Y3_N3
\Mux92~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux92~9_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux92~22_combout\))))) # (\R.curInst\(22) & (((!\Mux92~22_combout\ & ((\RegFile[28][30]~q\))) # (\Mux92~22_combout\ & (\RegFile[29][30]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux92~22_combout\)))) # (\R.curInst\(22) & ((!\Mux92~22_combout\ & (\RegFile[30][30]~q\)) # (\Mux92~22_combout\ & ((\RegFile[31][30]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[29][30]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[30][30]~q\,
	datad => \ALT_INV_RegFile[31][30]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux92~22_combout\,
	datag => \ALT_INV_RegFile[28][30]~q\,
	combout => \Mux92~9_combout\);

-- Location: FF_X62_Y5_N56
\RegFile[21][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(30),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][30]~q\);

-- Location: MLABCELL_X59_Y1_N48
\RegFile[22][30]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[22][30]~feeder_combout\ = ( \R.regWriteData\(30) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(30),
	combout => \RegFile[22][30]~feeder_combout\);

-- Location: FF_X59_Y1_N49
\RegFile[22][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[22][30]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][30]~q\);

-- Location: FF_X64_Y1_N56
\RegFile[17][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(30),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][30]~q\);

-- Location: MLABCELL_X59_Y3_N39
\RegFile[18][30]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[18][30]~feeder_combout\ = ( \R.regWriteData\(30) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(30),
	combout => \RegFile[18][30]~feeder_combout\);

-- Location: FF_X59_Y3_N40
\RegFile[18][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][30]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][30]~q\);

-- Location: FF_X64_Y2_N50
\RegFile[19][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(30),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][30]~q\);

-- Location: LABCELL_X64_Y1_N3
\RegFile[16][30]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[16][30]~feeder_combout\ = \R.regWriteData\(30)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101010101010101010101010101010101010101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.regWriteData\(30),
	combout => \RegFile[16][30]~feeder_combout\);

-- Location: FF_X64_Y1_N5
\RegFile[16][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[16][30]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][30]~q\);

-- Location: LABCELL_X64_Y1_N54
\Mux92~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux92~18_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[16][30]~q\))) # (\R.curInst\(20) & (\RegFile[17][30]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & (\RegFile[18][30]~q\)) # (\R.curInst\(20) & ((\RegFile[19][30]~q\)))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001110111011101110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[17][30]~q\,
	datac => \ALT_INV_RegFile[18][30]~q\,
	datad => \ALT_INV_RegFile[19][30]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][30]~q\,
	combout => \Mux92~18_combout\);

-- Location: MLABCELL_X59_Y3_N57
\RegFile[20][30]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[20][30]~feeder_combout\ = ( \R.regWriteData\(30) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(30),
	combout => \RegFile[20][30]~feeder_combout\);

-- Location: FF_X59_Y3_N58
\RegFile[20][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[20][30]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][30]~q\);

-- Location: LABCELL_X62_Y5_N18
\Mux92~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux92~5_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux92~18_combout\))))) # (\R.curInst\(22) & (((!\Mux92~18_combout\ & ((\RegFile[20][30]~q\))) # (\Mux92~18_combout\ & (\RegFile[21][30]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux92~18_combout\)))) # (\R.curInst\(22) & ((!\Mux92~18_combout\ & (\RegFile[22][30]~q\)) # (\Mux92~18_combout\ & ((\RegFile[23][30]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][30]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[22][30]~q\,
	datad => \ALT_INV_RegFile[23][30]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux92~18_combout\,
	datag => \ALT_INV_RegFile[20][30]~q\,
	combout => \Mux92~5_combout\);

-- Location: FF_X67_Y3_N38
\RegFile[3][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(30),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][30]~q\);

-- Location: FF_X61_Y5_N38
\RegFile[2][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(30),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][30]~q\);

-- Location: FF_X67_Y3_N29
\RegFile[6][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(30),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][30]~q\);

-- Location: FF_X67_Y5_N7
\RegFile[4][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(30),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][30]~q\);

-- Location: FF_X67_Y3_N55
\RegFile[7][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(30),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][30]~q\);

-- Location: FF_X62_Y3_N58
\RegFile[5][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(30),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][30]~q\);

-- Location: LABCELL_X62_Y3_N57
\Mux92~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux92~0_combout\ = ( \RegFile[5][30]~q\ & ( \R.curInst\(21) & ( (!\R.curInst\(20) & (\RegFile[6][30]~q\)) # (\R.curInst\(20) & ((\RegFile[7][30]~q\))) ) ) ) # ( !\RegFile[5][30]~q\ & ( \R.curInst\(21) & ( (!\R.curInst\(20) & (\RegFile[6][30]~q\)) # 
-- (\R.curInst\(20) & ((\RegFile[7][30]~q\))) ) ) ) # ( \RegFile[5][30]~q\ & ( !\R.curInst\(21) & ( (\R.curInst\(20)) # (\RegFile[4][30]~q\) ) ) ) # ( !\RegFile[5][30]~q\ & ( !\R.curInst\(21) & ( (\RegFile[4][30]~q\ & !\R.curInst\(20)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100000000001100111111111101010101000011110101010100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[6][30]~q\,
	datab => \ALT_INV_RegFile[4][30]~q\,
	datac => \ALT_INV_RegFile[7][30]~q\,
	datad => \ALT_INV_R.curInst\(20),
	datae => \ALT_INV_RegFile[5][30]~q\,
	dataf => \ALT_INV_R.curInst\(21),
	combout => \Mux92~0_combout\);

-- Location: LABCELL_X61_Y5_N12
\RegFile[1][30]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[1][30]~feeder_combout\ = \R.regWriteData\(30)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.regWriteData\(30),
	combout => \RegFile[1][30]~feeder_combout\);

-- Location: FF_X61_Y5_N14
\RegFile[1][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[1][30]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][30]~q\);

-- Location: LABCELL_X61_Y5_N36
\Mux92~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux92~26_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((\RegFile[1][30]~q\ & (\R.curInst\(20)))))) # (\R.curInst\(22) & ((((\Mux92~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (((\RegFile[2][30]~q\)))) # 
-- (\R.curInst\(20) & (\RegFile[3][30]~q\)))) # (\R.curInst\(22) & ((((\Mux92~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001010000010100010001001010101010111110101111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[3][30]~q\,
	datac => \ALT_INV_RegFile[2][30]~q\,
	datad => \ALT_INV_R.curInst\(20),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux92~0_combout\,
	datag => \ALT_INV_RegFile[1][30]~q\,
	combout => \Mux92~26_combout\);

-- Location: FF_X62_Y2_N50
\RegFile[13][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(30),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][30]~q\);

-- Location: FF_X70_Y2_N56
\RegFile[15][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(30),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][30]~q\);

-- Location: FF_X62_Y2_N20
\RegFile[14][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(30),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][30]~q\);

-- Location: FF_X70_Y2_N14
\RegFile[11][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(30),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][30]~q\);

-- Location: FF_X70_Y2_N32
\RegFile[9][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(30),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][30]~q\);

-- Location: MLABCELL_X59_Y3_N30
\RegFile[10][30]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[10][30]~feeder_combout\ = ( \R.regWriteData\(30) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(30),
	combout => \RegFile[10][30]~feeder_combout\);

-- Location: FF_X59_Y3_N32
\RegFile[10][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[10][30]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][30]~q\);

-- Location: MLABCELL_X59_Y1_N9
\RegFile[8][30]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[8][30]~feeder_combout\ = ( \R.regWriteData\(30) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(30),
	combout => \RegFile[8][30]~feeder_combout\);

-- Location: FF_X59_Y1_N10
\RegFile[8][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[8][30]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][30]~q\);

-- Location: LABCELL_X70_Y2_N30
\Mux92~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux92~14_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[8][30]~q\))) # (\R.curInst\(20) & (\RegFile[9][30]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[10][30]~q\))) # (\R.curInst\(20) & (\RegFile[11][30]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[11][30]~q\,
	datab => \ALT_INV_RegFile[9][30]~q\,
	datac => \ALT_INV_RegFile[10][30]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][30]~q\,
	combout => \Mux92~14_combout\);

-- Location: FF_X62_Y2_N26
\RegFile[12][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(30),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][30]~q\);

-- Location: LABCELL_X67_Y2_N42
\Mux92~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux92~1_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux92~14_combout\)))) # (\R.curInst\(22) & ((!\Mux92~14_combout\ & ((\RegFile[12][30]~q\))) # (\Mux92~14_combout\ & (\RegFile[13][30]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux92~14_combout\)))) # (\R.curInst\(22) & ((!\Mux92~14_combout\ & ((\RegFile[14][30]~q\))) # (\Mux92~14_combout\ & (\RegFile[15][30]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][30]~q\,
	datab => \ALT_INV_RegFile[15][30]~q\,
	datac => \ALT_INV_RegFile[14][30]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux92~14_combout\,
	datag => \ALT_INV_RegFile[12][30]~q\,
	combout => \Mux92~1_combout\);

-- Location: LABCELL_X61_Y5_N51
\Mux92~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux92~13_combout\ = ( \Mux92~26_combout\ & ( \Mux92~1_combout\ & ( (!\R.curInst\(24)) # ((!\R.curInst\(23) & ((\Mux92~5_combout\))) # (\R.curInst\(23) & (\Mux92~9_combout\))) ) ) ) # ( !\Mux92~26_combout\ & ( \Mux92~1_combout\ & ( (!\R.curInst\(23) & 
-- (((\Mux92~5_combout\ & \R.curInst\(24))))) # (\R.curInst\(23) & (((!\R.curInst\(24))) # (\Mux92~9_combout\))) ) ) ) # ( \Mux92~26_combout\ & ( !\Mux92~1_combout\ & ( (!\R.curInst\(23) & (((!\R.curInst\(24)) # (\Mux92~5_combout\)))) # (\R.curInst\(23) & 
-- (\Mux92~9_combout\ & ((\R.curInst\(24))))) ) ) ) # ( !\Mux92~26_combout\ & ( !\Mux92~1_combout\ & ( (\R.curInst\(24) & ((!\R.curInst\(23) & ((\Mux92~5_combout\))) # (\R.curInst\(23) & (\Mux92~9_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000011011101010100001101101010101000110111111111100011011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(23),
	datab => \ALT_INV_Mux92~9_combout\,
	datac => \ALT_INV_Mux92~5_combout\,
	datad => \ALT_INV_R.curInst\(24),
	datae => \ALT_INV_Mux92~26_combout\,
	dataf => \ALT_INV_Mux92~1_combout\,
	combout => \Mux92~13_combout\);

-- Location: LABCELL_X60_Y5_N54
\NxR.aluData2[30]~30\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[30]~30_combout\ = ( \Mux124~1_combout\ & ( \Mux92~13_combout\ & ( (!\vAluSrc2~1_combout\) # (\Equal4~1_combout\) ) ) ) # ( !\Mux124~1_combout\ & ( \Mux92~13_combout\ & ( !\vAluSrc2~1_combout\ ) ) ) # ( \Mux124~1_combout\ & ( 
-- !\Mux92~13_combout\ & ( (\Equal4~1_combout\ & \vAluSrc2~1_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000110000001111110000111100001111001111110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Equal4~1_combout\,
	datac => \ALT_INV_vAluSrc2~1_combout\,
	datae => \ALT_INV_Mux124~1_combout\,
	dataf => \ALT_INV_Mux92~13_combout\,
	combout => \NxR.aluData2[30]~30_combout\);

-- Location: FF_X60_Y5_N55
\R.aluData2[30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR.aluData2[30]~30_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData2\(30));

-- Location: FF_X73_Y5_N22
\R.aluData1[30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux224~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData1\(30));

-- Location: MLABCELL_X78_Y5_N27
\Add1~117\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~117_sumout\ = SUM(( \R.aluData1\(29) ) + ( \R.aluData2\(29) ) + ( \Add1~114\ ))
-- \Add1~118\ = CARRY(( \R.aluData1\(29) ) + ( \R.aluData2\(29) ) + ( \Add1~114\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData1\(29),
	dataf => \ALT_INV_R.aluData2\(29),
	cin => \Add1~114\,
	sumout => \Add1~117_sumout\,
	cout => \Add1~118\);

-- Location: MLABCELL_X78_Y5_N30
\Add1~121\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~121_sumout\ = SUM(( \R.aluData1\(30) ) + ( \R.aluData2\(30) ) + ( \Add1~118\ ))
-- \Add1~122\ = CARRY(( \R.aluData1\(30) ) + ( \R.aluData2\(30) ) + ( \Add1~118\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluData2\(30),
	datad => \ALT_INV_R.aluData1\(30),
	cin => \Add1~118\,
	sumout => \Add1~121_sumout\,
	cout => \Add1~122\);

-- Location: LABCELL_X75_Y4_N6
\Mux129~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux129~0_combout\ = ( \R.curInst\(25) & ( ((\vAluSrc1~0_combout\ & ((\Mux124~0_combout\) # (\R.curInst\(2))))) # (\Mux123~1_combout\) ) ) # ( !\R.curInst\(25) & ( ((\vAluSrc1~0_combout\ & \Mux124~0_combout\)) # (\Mux123~1_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010111111111000001011111111100010101111111110001010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluSrc1~0_combout\,
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_Mux124~0_combout\,
	datad => \ALT_INV_Mux123~1_combout\,
	dataf => \ALT_INV_R.curInst\(25),
	combout => \Mux129~0_combout\);

-- Location: FF_X62_Y1_N41
\RegFile[2][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(25),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][25]~q\);

-- Location: FF_X68_Y3_N2
\RegFile[3][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(25),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][25]~q\);

-- Location: FF_X59_Y5_N49
\RegFile[6][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(25),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][25]~q\);

-- Location: FF_X68_Y3_N13
\RegFile[7][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(25),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][25]~q\);

-- Location: LABCELL_X60_Y3_N0
\RegFile[4][25]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[4][25]~feeder_combout\ = ( \R.regWriteData\(25) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(25),
	combout => \RegFile[4][25]~feeder_combout\);

-- Location: FF_X60_Y3_N1
\RegFile[4][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[4][25]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][25]~q\);

-- Location: LABCELL_X60_Y3_N21
\RegFile[5][25]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[5][25]~feeder_combout\ = ( \R.regWriteData\(25) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(25),
	combout => \RegFile[5][25]~feeder_combout\);

-- Location: FF_X60_Y3_N22
\RegFile[5][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[5][25]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][25]~q\);

-- Location: LABCELL_X61_Y1_N51
\Mux97~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux97~0_combout\ = ( \R.curInst\(20) & ( \R.curInst\(21) & ( \RegFile[7][25]~q\ ) ) ) # ( !\R.curInst\(20) & ( \R.curInst\(21) & ( \RegFile[6][25]~q\ ) ) ) # ( \R.curInst\(20) & ( !\R.curInst\(21) & ( \RegFile[5][25]~q\ ) ) ) # ( !\R.curInst\(20) & ( 
-- !\R.curInst\(21) & ( \RegFile[4][25]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000000001111111101010101010101010011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[6][25]~q\,
	datab => \ALT_INV_RegFile[7][25]~q\,
	datac => \ALT_INV_RegFile[4][25]~q\,
	datad => \ALT_INV_RegFile[5][25]~q\,
	datae => \ALT_INV_R.curInst\(20),
	dataf => \ALT_INV_R.curInst\(21),
	combout => \Mux97~0_combout\);

-- Location: FF_X61_Y5_N17
\RegFile[1][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(25),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][25]~q\);

-- Location: LABCELL_X62_Y1_N39
\Mux97~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux97~26_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (\R.curInst\(20) & (\RegFile[1][25]~q\))) # (\R.curInst\(22) & ((((\Mux97~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (\RegFile[2][25]~q\)) # 
-- (\R.curInst\(20) & (((\RegFile[3][25]~q\)))))) # (\R.curInst\(22) & ((((\Mux97~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010000000100000010000100110000110111001101110011101101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(20),
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[2][25]~q\,
	datad => \ALT_INV_RegFile[3][25]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux97~0_combout\,
	datag => \ALT_INV_RegFile[1][25]~q\,
	combout => \Mux97~26_combout\);

-- Location: LABCELL_X68_Y1_N48
\RegFile[30][25]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[30][25]~feeder_combout\ = ( \R.regWriteData\(25) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(25),
	combout => \RegFile[30][25]~feeder_combout\);

-- Location: FF_X68_Y1_N49
\RegFile[30][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[30][25]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][25]~q\);

-- Location: FF_X62_Y1_N14
\RegFile[29][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(25),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][25]~q\);

-- Location: FF_X67_Y1_N20
\RegFile[25][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(25),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][25]~q\);

-- Location: FF_X67_Y2_N35
\RegFile[26][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(25),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][25]~q\);

-- Location: FF_X67_Y1_N50
\RegFile[27][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(25),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][25]~q\);

-- Location: MLABCELL_X59_Y2_N57
\RegFile[24][25]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[24][25]~feeder_combout\ = ( \R.regWriteData\(25) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(25),
	combout => \RegFile[24][25]~feeder_combout\);

-- Location: FF_X59_Y2_N58
\RegFile[24][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[24][25]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][25]~q\);

-- Location: LABCELL_X67_Y1_N18
\Mux97~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux97~22_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[24][25]~q\))) # (\R.curInst\(20) & (\RegFile[25][25]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & (\RegFile[26][25]~q\)) # (\R.curInst\(20) & ((\RegFile[27][25]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[25][25]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[26][25]~q\,
	datad => \ALT_INV_RegFile[27][25]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][25]~q\,
	combout => \Mux97~22_combout\);

-- Location: LABCELL_X73_Y2_N0
\RegFile[28][25]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[28][25]~feeder_combout\ = ( \R.regWriteData\(25) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(25),
	combout => \RegFile[28][25]~feeder_combout\);

-- Location: FF_X73_Y2_N1
\RegFile[28][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[28][25]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][25]~q\);

-- Location: LABCELL_X62_Y1_N12
\Mux97~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux97~9_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux97~22_combout\)))) # (\R.curInst\(22) & ((!\Mux97~22_combout\ & (\RegFile[28][25]~q\)) # (\Mux97~22_combout\ & ((\RegFile[29][25]~q\)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) 
-- & ((((\Mux97~22_combout\))))) # (\R.curInst\(22) & (((!\Mux97~22_combout\ & ((\RegFile[30][25]~q\))) # (\Mux97~22_combout\ & (\RegFile[31][25]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111001100111111111101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][25]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[30][25]~q\,
	datad => \ALT_INV_RegFile[29][25]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux97~22_combout\,
	datag => \ALT_INV_RegFile[28][25]~q\,
	combout => \Mux97~9_combout\);

-- Location: FF_X68_Y2_N50
\RegFile[15][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(25),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][25]~q\);

-- Location: FF_X62_Y2_N14
\RegFile[13][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(25),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][25]~q\);

-- Location: LABCELL_X62_Y2_N21
\RegFile[14][25]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[14][25]~feeder_combout\ = ( \R.regWriteData\(25) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(25),
	combout => \RegFile[14][25]~feeder_combout\);

-- Location: FF_X62_Y2_N22
\RegFile[14][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[14][25]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][25]~q\);

-- Location: FF_X68_Y2_N38
\RegFile[11][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(25),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][25]~q\);

-- Location: FF_X68_Y2_N8
\RegFile[9][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(25),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][25]~q\);

-- Location: FF_X64_Y3_N49
\RegFile[10][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(25),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][25]~q\);

-- Location: FF_X63_Y6_N22
\RegFile[8][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(25),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][25]~q\);

-- Location: LABCELL_X68_Y2_N6
\Mux97~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux97~14_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[8][25]~q\))) # (\R.curInst\(20) & (\RegFile[9][25]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[10][25]~q\))) # (\R.curInst\(20) & (\RegFile[11][25]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[11][25]~q\,
	datab => \ALT_INV_RegFile[9][25]~q\,
	datac => \ALT_INV_RegFile[10][25]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][25]~q\,
	combout => \Mux97~14_combout\);

-- Location: LABCELL_X62_Y2_N27
\RegFile[12][25]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[12][25]~feeder_combout\ = ( \R.regWriteData\(25) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(25),
	combout => \RegFile[12][25]~feeder_combout\);

-- Location: FF_X62_Y2_N29
\RegFile[12][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[12][25]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][25]~q\);

-- Location: LABCELL_X62_Y2_N12
\Mux97~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux97~1_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux97~14_combout\)))) # (\R.curInst\(22) & ((!\Mux97~14_combout\ & ((\RegFile[12][25]~q\))) # (\Mux97~14_combout\ & (\RegFile[13][25]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux97~14_combout\)))) # (\R.curInst\(22) & ((!\Mux97~14_combout\ & ((\RegFile[14][25]~q\))) # (\Mux97~14_combout\ & (\RegFile[15][25]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][25]~q\,
	datab => \ALT_INV_RegFile[13][25]~q\,
	datac => \ALT_INV_RegFile[14][25]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux97~14_combout\,
	datag => \ALT_INV_RegFile[12][25]~q\,
	combout => \Mux97~1_combout\);

-- Location: FF_X61_Y6_N55
\RegFile[21][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(25),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][25]~q\);

-- Location: FF_X61_Y6_N25
\RegFile[22][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(25),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][25]~q\);

-- Location: FF_X64_Y2_N8
\RegFile[23][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(25),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][25]~q\);

-- Location: FF_X64_Y2_N2
\RegFile[17][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(25),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][25]~q\);

-- Location: FF_X64_Y2_N14
\RegFile[19][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(25),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][25]~q\);

-- Location: MLABCELL_X59_Y3_N42
\RegFile[18][25]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[18][25]~feeder_combout\ = ( \R.regWriteData\(25) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(25),
	combout => \RegFile[18][25]~feeder_combout\);

-- Location: FF_X59_Y3_N43
\RegFile[18][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][25]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][25]~q\);

-- Location: LABCELL_X64_Y1_N30
\RegFile[16][25]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[16][25]~feeder_combout\ = ( \R.regWriteData\(25) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(25),
	combout => \RegFile[16][25]~feeder_combout\);

-- Location: FF_X64_Y1_N31
\RegFile[16][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[16][25]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][25]~q\);

-- Location: LABCELL_X64_Y2_N0
\Mux97~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux97~18_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[16][25]~q\))) # (\R.curInst\(20) & (\RegFile[17][25]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[18][25]~q\))) # (\R.curInst\(20) & (\RegFile[19][25]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[17][25]~q\,
	datab => \ALT_INV_RegFile[19][25]~q\,
	datac => \ALT_INV_RegFile[18][25]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][25]~q\,
	combout => \Mux97~18_combout\);

-- Location: MLABCELL_X59_Y3_N18
\RegFile[20][25]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[20][25]~feeder_combout\ = ( \R.regWriteData\(25) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(25),
	combout => \RegFile[20][25]~feeder_combout\);

-- Location: FF_X59_Y3_N19
\RegFile[20][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[20][25]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][25]~q\);

-- Location: LABCELL_X62_Y2_N54
\Mux97~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux97~5_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux97~18_combout\))))) # (\R.curInst\(22) & (((!\Mux97~18_combout\ & ((\RegFile[20][25]~q\))) # (\Mux97~18_combout\ & (\RegFile[21][25]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux97~18_combout\)))) # (\R.curInst\(22) & ((!\Mux97~18_combout\ & (\RegFile[22][25]~q\)) # (\Mux97~18_combout\ & ((\RegFile[23][25]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][25]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[22][25]~q\,
	datad => \ALT_INV_RegFile[23][25]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux97~18_combout\,
	datag => \ALT_INV_RegFile[20][25]~q\,
	combout => \Mux97~5_combout\);

-- Location: LABCELL_X62_Y1_N45
\Mux97~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux97~13_combout\ = ( \Mux97~1_combout\ & ( \Mux97~5_combout\ & ( (!\R.curInst\(23) & (((\R.curInst\(24))) # (\Mux97~26_combout\))) # (\R.curInst\(23) & (((!\R.curInst\(24)) # (\Mux97~9_combout\)))) ) ) ) # ( !\Mux97~1_combout\ & ( \Mux97~5_combout\ & ( 
-- (!\R.curInst\(23) & (((\R.curInst\(24))) # (\Mux97~26_combout\))) # (\R.curInst\(23) & (((\Mux97~9_combout\ & \R.curInst\(24))))) ) ) ) # ( \Mux97~1_combout\ & ( !\Mux97~5_combout\ & ( (!\R.curInst\(23) & (\Mux97~26_combout\ & ((!\R.curInst\(24))))) # 
-- (\R.curInst\(23) & (((!\R.curInst\(24)) # (\Mux97~9_combout\)))) ) ) ) # ( !\Mux97~1_combout\ & ( !\Mux97~5_combout\ & ( (!\R.curInst\(23) & (\Mux97~26_combout\ & ((!\R.curInst\(24))))) # (\R.curInst\(23) & (((\Mux97~9_combout\ & \R.curInst\(24))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010001000000101011101110000010100100010101011110111011110101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(23),
	datab => \ALT_INV_Mux97~26_combout\,
	datac => \ALT_INV_Mux97~9_combout\,
	datad => \ALT_INV_R.curInst\(24),
	datae => \ALT_INV_Mux97~1_combout\,
	dataf => \ALT_INV_Mux97~5_combout\,
	combout => \Mux97~13_combout\);

-- Location: LABCELL_X79_Y5_N54
\NxR.aluData2[25]~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[25]~22_combout\ = ( \Mux97~13_combout\ & ( (!\vAluSrc2~1_combout\) # ((\Mux129~0_combout\ & \Equal4~1_combout\)) ) ) # ( !\Mux97~13_combout\ & ( (\Mux129~0_combout\ & (\vAluSrc2~1_combout\ & \Equal4~1_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000011000000000000001111110000111100111111000011110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Mux129~0_combout\,
	datac => \ALT_INV_vAluSrc2~1_combout\,
	datad => \ALT_INV_Equal4~1_combout\,
	dataf => \ALT_INV_Mux97~13_combout\,
	combout => \NxR.aluData2[25]~22_combout\);

-- Location: FF_X79_Y5_N56
\R.aluData2[25]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR.aluData2[25]~22_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData2[25]~DUPLICATE_q\);

-- Location: FF_X74_Y3_N58
\R.aluData1[24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux230~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData1\(24));

-- Location: FF_X74_Y5_N28
\R.aluData1[21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux233~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData1\(21));

-- Location: LABCELL_X74_Y4_N21
\Mux134~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux134~0_combout\ = ( \R.curInst\(20) & ( ((\vAluSrc1~0_combout\ & ((\Mux124~0_combout\) # (\R.curInst\(2))))) # (\Mux123~1_combout\) ) ) # ( !\R.curInst\(20) & ( ((\vAluSrc1~0_combout\ & \Mux124~0_combout\)) # (\Mux123~1_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111101011111000011110101111100011111010111110001111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluSrc1~0_combout\,
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_Mux123~1_combout\,
	datad => \ALT_INV_Mux124~0_combout\,
	dataf => \ALT_INV_R.curInst\(20),
	combout => \Mux134~0_combout\);

-- Location: LABCELL_X81_Y6_N54
\Add0~73\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~73_sumout\ = SUM(( \R.curPC\(20) ) + ( GND ) + ( \Add0~70\ ))
-- \Add0~74\ = CARRY(( \R.curPC\(20) ) + ( GND ) + ( \Add0~70\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.curPC\(20),
	cin => \Add0~70\,
	sumout => \Add0~73_sumout\,
	cout => \Add0~74\);

-- Location: LABCELL_X79_Y8_N12
\R.regWriteData[20]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.regWriteData[20]~feeder_combout\ = ( \Add0~73_sumout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_Add0~73_sumout\,
	combout => \R.regWriteData[20]~feeder_combout\);

-- Location: LABCELL_X71_Y7_N12
\ShiftRight0~7_RTM0235\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight0~7_RTM0235_combout\ = ( \Mux151~0_combout\ & ( \Mux119~13_combout\ & ( (!\vAluSrc2~1_combout\) # (\Equal4~1_combout\) ) ) ) # ( !\Mux151~0_combout\ & ( \Mux119~13_combout\ & ( (!\vAluSrc2~1_combout\) # ((\Equal4~1_combout\ & 
-- \Mux152~0_combout\)) ) ) ) # ( \Mux151~0_combout\ & ( !\Mux119~13_combout\ & ( (!\vAluSrc2~1_combout\ & (\Mux120~13_combout\)) # (\vAluSrc2~1_combout\ & ((\Equal4~1_combout\))) ) ) ) # ( !\Mux151~0_combout\ & ( !\Mux119~13_combout\ & ( 
-- (!\vAluSrc2~1_combout\ & (\Mux120~13_combout\)) # (\vAluSrc2~1_combout\ & (((\Equal4~1_combout\ & \Mux152~0_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100010001000111010001110100011111001100110011111100111111001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux120~13_combout\,
	datab => \ALT_INV_vAluSrc2~1_combout\,
	datac => \ALT_INV_Equal4~1_combout\,
	datad => \ALT_INV_Mux152~0_combout\,
	datae => \ALT_INV_Mux151~0_combout\,
	dataf => \ALT_INV_Mux119~13_combout\,
	combout => \ShiftRight0~7_RTM0235_combout\);

-- Location: FF_X71_Y7_N13
\ShiftRight0~7_OTERM233DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight0~7_RTM0235_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight0~7_OTERM233DUPLICATE_q\);

-- Location: LABCELL_X71_Y7_N30
\ShiftLeft0~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~4_combout\ = ( !\NxR.aluData2[1]~17_combout\ & ( (\NxR.aluData2[2]~19_combout\ & (!\NxR.aluData2[0]~16_combout\ & (\Mux254~0_combout\ & !\NxR.aluData2[3]~18_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010000000000000001000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_NxR.aluData2[2]~19_combout\,
	datab => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datac => \ALT_INV_Mux254~0_combout\,
	datad => \ALT_INV_NxR.aluData2[3]~18_combout\,
	dataf => \ALT_INV_NxR.aluData2[1]~17_combout\,
	combout => \ShiftLeft0~4_combout\);

-- Location: FF_X71_Y7_N31
\ShiftLeft0~4_NEW_REG236\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~4_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~4_OTERM237\);

-- Location: FF_X73_Y5_N10
\R.aluData1[20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux234~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData1\(20));

-- Location: MLABCELL_X84_Y5_N18
\Selector12~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector12~3_combout\ = ( \R.aluData1\(20) & ( \R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( (!\R.aluOp.ALUOpOr~q\ & (!\R.aluOp.ALUOpXor~DUPLICATE_q\ & !\R.aluData2\(20))) ) ) ) # ( !\R.aluData1\(20) & ( \R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( (!\R.aluData2\(20)) # 
-- ((!\R.aluOp.ALUOpOr~q\ & !\R.aluOp.ALUOpXor~DUPLICATE_q\)) ) ) ) # ( \R.aluData1\(20) & ( !\R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( (!\R.aluOp.ALUOpOr~q\ & ((!\R.aluOp.ALUOpXor~DUPLICATE_q\) # (\R.aluData2\(20)))) ) ) ) # ( !\R.aluData1\(20) & ( 
-- !\R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( (!\R.aluData2\(20)) # ((!\R.aluOp.ALUOpOr~q\ & !\R.aluOp.ALUOpXor~DUPLICATE_q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111100011111000100010101000101011111000111110001000000010000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpOr~q\,
	datab => \ALT_INV_R.aluOp.ALUOpXor~DUPLICATE_q\,
	datac => \ALT_INV_R.aluData2\(20),
	datae => \ALT_INV_R.aluData1\(20),
	dataf => \ALT_INV_R.aluOp.ALUOpAnd~DUPLICATE_q\,
	combout => \Selector12~3_combout\);

-- Location: LABCELL_X81_Y7_N18
\Selector12~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector12~4_combout\ = ( \ShiftLeft0~4_OTERM237\ & ( \Selector12~3_combout\ & ( (!\Selector12~2_OTERM395\ & !\Selector17~0_OTERM391\) ) ) ) # ( !\ShiftLeft0~4_OTERM237\ & ( \Selector12~3_combout\ & ( (!\Selector17~0_OTERM391\ & 
-- ((!\Selector12~2_OTERM395\) # ((!\ShiftLeft0~5_OTERM203\) # (\ShiftRight0~7_OTERM233DUPLICATE_q\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011110000101100001010000010100000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector12~2_OTERM395\,
	datab => \ALT_INV_ShiftRight0~7_OTERM233DUPLICATE_q\,
	datac => \ALT_INV_Selector17~0_OTERM391\,
	datad => \ALT_INV_ShiftLeft0~5_OTERM203\,
	datae => \ALT_INV_ShiftLeft0~4_OTERM237\,
	dataf => \ALT_INV_Selector12~3_combout\,
	combout => \Selector12~4_combout\);

-- Location: MLABCELL_X78_Y8_N12
\Comb:vRegWriteData[20]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[20]~3_combout\ = ( \R.memToReg~q\ & ( (\Selector12~4_combout\ & (!\Selector12~1_combout\ & \R.aluCalc~q\)) ) ) # ( !\R.memToReg~q\ & ( (!\R.aluCalc~q\ & (!\R.aluRes\(20))) # (\R.aluCalc~q\ & (((\Selector12~4_combout\ & 
-- !\Selector12~1_combout\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010101000110000101010100011000000000000001100000000000000110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluRes\(20),
	datab => \ALT_INV_Selector12~4_combout\,
	datac => \ALT_INV_Selector12~1_combout\,
	datad => \ALT_INV_R.aluCalc~q\,
	dataf => \ALT_INV_R.memToReg~q\,
	combout => \Comb:vRegWriteData[20]~3_combout\);

-- Location: LABCELL_X75_Y4_N48
\Mux137~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux137~0_combout\ = ( \Mux123~2_combout\ & ( \R.curInst\(17) ) ) # ( !\Mux123~2_combout\ & ( \R.curInst\(17) & ( ((\vAluSrc1~0_combout\ & ((\R.curInst\(2)) # (\Mux124~0_combout\)))) # (\Mux149~0_combout\) ) ) ) # ( \Mux123~2_combout\ & ( !\R.curInst\(17) 
-- ) ) # ( !\Mux123~2_combout\ & ( !\R.curInst\(17) & ( (\Mux124~0_combout\ & \vAluSrc1~0_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010101111111111111111100001111011111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux124~0_combout\,
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_Mux149~0_combout\,
	datad => \ALT_INV_vAluSrc1~0_combout\,
	datae => \ALT_INV_Mux123~2_combout\,
	dataf => \ALT_INV_R.curInst\(17),
	combout => \Mux137~0_combout\);

-- Location: LABCELL_X75_Y4_N57
\Mux139~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux139~0_combout\ = ( \Mux123~2_combout\ & ( \R.curInst\(15) ) ) # ( !\Mux123~2_combout\ & ( \R.curInst\(15) & ( ((\vAluSrc1~0_combout\ & ((\R.curInst\(2)) # (\Mux124~0_combout\)))) # (\Mux149~0_combout\) ) ) ) # ( \Mux123~2_combout\ & ( !\R.curInst\(15) 
-- ) ) # ( !\Mux123~2_combout\ & ( !\R.curInst\(15) & ( (\Mux124~0_combout\ & \vAluSrc1~0_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101111111111111111100000111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux124~0_combout\,
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_vAluSrc1~0_combout\,
	datad => \ALT_INV_Mux149~0_combout\,
	datae => \ALT_INV_Mux123~2_combout\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux139~0_combout\);

-- Location: LABCELL_X81_Y6_N33
\Add0~45\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~45_sumout\ = SUM(( \R.curPC\(13) ) + ( GND ) + ( \Add0~42\ ))
-- \Add0~46\ = CARRY(( \R.curPC\(13) ) + ( GND ) + ( \Add0~42\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.curPC\(13),
	cin => \Add0~42\,
	sumout => \Add0~45_sumout\,
	cout => \Add0~46\);

-- Location: LABCELL_X81_Y6_N36
\Add0~49\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~49_sumout\ = SUM(( \R.curPC\(14) ) + ( GND ) + ( \Add0~46\ ))
-- \Add0~50\ = CARRY(( \R.curPC\(14) ) + ( GND ) + ( \Add0~46\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.curPC\(14),
	cin => \Add0~46\,
	sumout => \Add0~49_sumout\,
	cout => \Add0~50\);

-- Location: LABCELL_X81_Y6_N39
\Add0~53\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~53_sumout\ = SUM(( \R.curPC\(15) ) + ( GND ) + ( \Add0~50\ ))
-- \Add0~54\ = CARRY(( \R.curPC\(15) ) + ( GND ) + ( \Add0~50\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curPC\(15),
	cin => \Add0~50\,
	sumout => \Add0~53_sumout\,
	cout => \Add0~54\);

-- Location: LABCELL_X80_Y6_N24
\R.regWriteData[15]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.regWriteData[15]~feeder_combout\ = \Add0~53_sumout\

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Add0~53_sumout\,
	combout => \R.regWriteData[15]~feeder_combout\);

-- Location: FF_X74_Y2_N26
\RegFile[29][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(15),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][15]~q\);

-- Location: FF_X75_Y2_N16
\RegFile[30][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(15),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][15]~q\);

-- Location: FF_X67_Y2_N55
\RegFile[27][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(15),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][15]~q\);

-- Location: FF_X67_Y2_N32
\RegFile[26][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(15),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][15]~q\);

-- Location: FF_X67_Y2_N14
\RegFile[25][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(15),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][15]~q\);

-- Location: FF_X59_Y2_N16
\RegFile[24][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(15),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][15]~q\);

-- Location: MLABCELL_X72_Y2_N12
\Mux75~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux75~22_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & (\RegFile[24][15]~q\)) # (\R.curInst\(15) & ((\RegFile[25][15]~q\))))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & ((\RegFile[26][15]~q\))) # (\R.curInst\(15) & (\RegFile[27][15]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110000110011111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[27][15]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[26][15]~q\,
	datad => \ALT_INV_RegFile[25][15]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][15]~q\,
	combout => \Mux75~22_combout\);

-- Location: FF_X73_Y2_N43
\RegFile[28][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(15),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][15]~q\);

-- Location: MLABCELL_X72_Y2_N42
\Mux75~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux75~9_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux75~22_combout\)))) # (\R.curInst\(17) & ((!\Mux75~22_combout\ & ((\RegFile[28][15]~q\))) # (\Mux75~22_combout\ & (\RegFile[29][15]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux75~22_combout\)))) # (\R.curInst\(17) & ((!\Mux75~22_combout\ & ((\RegFile[30][15]~q\))) # (\Mux75~22_combout\ & (\RegFile[31][15]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][15]~q\,
	datab => \ALT_INV_RegFile[29][15]~q\,
	datac => \ALT_INV_RegFile[30][15]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux75~22_combout\,
	datag => \ALT_INV_RegFile[28][15]~q\,
	combout => \Mux75~9_combout\);

-- Location: FF_X72_Y2_N38
\RegFile[15][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(15),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][15]~q\);

-- Location: FF_X62_Y2_N37
\RegFile[14][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(15),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][15]~q\);

-- Location: FF_X74_Y2_N56
\RegFile[13][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(15),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][15]~q\);

-- Location: FF_X72_Y2_N11
\RegFile[11][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(15),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][15]~q\);

-- Location: FF_X75_Y2_N1
\RegFile[10][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(15),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][15]~q\);

-- Location: FF_X74_Y2_N8
\RegFile[9][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(15),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][15]~q\);

-- Location: FF_X68_Y5_N49
\RegFile[8][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(15),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][15]~q\);

-- Location: MLABCELL_X72_Y2_N9
\Mux75~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux75~14_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & (\RegFile[8][15]~q\)) # (\R.curInst\(15) & ((\RegFile[9][15]~q\))))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & ((\RegFile[10][15]~q\))) # (\R.curInst\(15) & (\RegFile[11][15]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110000110011111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[11][15]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[10][15]~q\,
	datad => \ALT_INV_RegFile[9][15]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][15]~q\,
	combout => \Mux75~14_combout\);

-- Location: LABCELL_X62_Y2_N24
\RegFile[12][15]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[12][15]~feeder_combout\ = \R.regWriteData\(15)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.regWriteData\(15),
	combout => \RegFile[12][15]~feeder_combout\);

-- Location: FF_X62_Y2_N25
\RegFile[12][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[12][15]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][15]~q\);

-- Location: MLABCELL_X72_Y2_N36
\Mux75~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux75~1_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux75~14_combout\))))) # (\R.curInst\(17) & (((!\Mux75~14_combout\ & (\RegFile[12][15]~q\)) # (\Mux75~14_combout\ & ((\RegFile[13][15]~q\)))))) ) ) # ( \R.curInst\(16) & ( 
-- (!\R.curInst\(17) & ((((\Mux75~14_combout\))))) # (\R.curInst\(17) & (((!\Mux75~14_combout\ & ((\RegFile[14][15]~q\))) # (\Mux75~14_combout\ & (\RegFile[15][15]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110101010111111111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[15][15]~q\,
	datac => \ALT_INV_RegFile[14][15]~q\,
	datad => \ALT_INV_RegFile[13][15]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux75~14_combout\,
	datag => \ALT_INV_RegFile[12][15]~q\,
	combout => \Mux75~1_combout\);

-- Location: FF_X73_Y3_N2
\RegFile[3][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(15),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][15]~q\);

-- Location: FF_X72_Y3_N50
\RegFile[2][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(15),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][15]~q\);

-- Location: LABCELL_X67_Y5_N57
\RegFile[4][15]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[4][15]~feeder_combout\ = ( \R.regWriteData\(15) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(15),
	combout => \RegFile[4][15]~feeder_combout\);

-- Location: FF_X67_Y5_N58
\RegFile[4][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[4][15]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][15]~q\);

-- Location: FF_X73_Y3_N38
\RegFile[6][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(15),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][15]~q\);

-- Location: FF_X72_Y4_N32
\RegFile[5][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(15),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][15]~q\);

-- Location: FF_X73_Y3_N31
\RegFile[7][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(15),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][15]~q\);

-- Location: LABCELL_X73_Y3_N30
\Mux75~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux75~0_combout\ = ( \RegFile[7][15]~q\ & ( \R.curInst\(15) & ( (\RegFile[5][15]~q\) # (\R.curInst\(16)) ) ) ) # ( !\RegFile[7][15]~q\ & ( \R.curInst\(15) & ( (!\R.curInst\(16) & \RegFile[5][15]~q\) ) ) ) # ( \RegFile[7][15]~q\ & ( !\R.curInst\(15) & ( 
-- (!\R.curInst\(16) & (\RegFile[4][15]~q\)) # (\R.curInst\(16) & ((\RegFile[6][15]~q\))) ) ) ) # ( !\RegFile[7][15]~q\ & ( !\R.curInst\(15) & ( (!\R.curInst\(16) & (\RegFile[4][15]~q\)) # (\R.curInst\(16) & ((\RegFile[6][15]~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010011100100111001001110010011100000000101010100101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(16),
	datab => \ALT_INV_RegFile[4][15]~q\,
	datac => \ALT_INV_RegFile[6][15]~q\,
	datad => \ALT_INV_RegFile[5][15]~q\,
	datae => \ALT_INV_RegFile[7][15]~q\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux75~0_combout\);

-- Location: FF_X72_Y3_N40
\RegFile[1][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(15),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][15]~q\);

-- Location: LABCELL_X73_Y3_N0
\Mux75~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux75~26_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (\RegFile[1][15]~q\ & (\R.curInst\(15)))) # (\R.curInst\(17) & (((\Mux75~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & ((!\R.curInst\(15) & (((\RegFile[2][15]~q\)))) # 
-- (\R.curInst\(15) & (\RegFile[3][15]~q\)))) # (\R.curInst\(17) & ((((\Mux75~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001100000011000100010000110011001111110011111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][15]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[2][15]~q\,
	datad => \ALT_INV_R.curInst\(15),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux75~0_combout\,
	datag => \ALT_INV_RegFile[1][15]~q\,
	combout => \Mux75~26_combout\);

-- Location: FF_X72_Y1_N56
\RegFile[23][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(15),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][15]~q\);

-- Location: LABCELL_X71_Y1_N24
\RegFile[22][15]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[22][15]~feeder_combout\ = \R.regWriteData\(15)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.regWriteData\(15),
	combout => \RegFile[22][15]~feeder_combout\);

-- Location: FF_X71_Y1_N25
\RegFile[22][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[22][15]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][15]~q\);

-- Location: FF_X71_Y1_N44
\RegFile[21][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(15),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][15]~q\);

-- Location: MLABCELL_X72_Y1_N42
\RegFile[17][15]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[17][15]~feeder_combout\ = ( \R.regWriteData\(15) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(15),
	combout => \RegFile[17][15]~feeder_combout\);

-- Location: FF_X72_Y1_N43
\RegFile[17][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[17][15]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][15]~q\);

-- Location: LABCELL_X73_Y1_N54
\RegFile[18][15]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[18][15]~feeder_combout\ = ( \R.regWriteData\(15) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(15),
	combout => \RegFile[18][15]~feeder_combout\);

-- Location: FF_X73_Y1_N56
\RegFile[18][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][15]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][15]~q\);

-- Location: FF_X73_Y1_N32
\RegFile[19][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(15),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][15]~q\);

-- Location: LABCELL_X74_Y1_N27
\RegFile[16][15]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[16][15]~feeder_combout\ = ( \R.regWriteData\(15) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(15),
	combout => \RegFile[16][15]~feeder_combout\);

-- Location: FF_X74_Y1_N29
\RegFile[16][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[16][15]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][15]~q\);

-- Location: LABCELL_X73_Y1_N30
\Mux75~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux75~18_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[16][15]~q\))) # (\R.curInst\(15) & (\RegFile[17][15]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & (\RegFile[18][15]~q\)) # (\R.curInst\(15) & ((\RegFile[19][15]~q\)))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001110111011101110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[17][15]~q\,
	datac => \ALT_INV_RegFile[18][15]~q\,
	datad => \ALT_INV_RegFile[19][15]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][15]~q\,
	combout => \Mux75~18_combout\);

-- Location: FF_X71_Y1_N49
\RegFile[20][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(15),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][15]~q\);

-- Location: MLABCELL_X72_Y1_N54
\Mux75~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux75~5_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux75~18_combout\)))) # (\R.curInst\(17) & ((!\Mux75~18_combout\ & (\RegFile[20][15]~q\)) # (\Mux75~18_combout\ & ((\RegFile[21][15]~q\)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) 
-- & ((((\Mux75~18_combout\))))) # (\R.curInst\(17) & (((!\Mux75~18_combout\ & ((\RegFile[22][15]~q\))) # (\Mux75~18_combout\ & (\RegFile[23][15]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111001100111111111101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[23][15]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[22][15]~q\,
	datad => \ALT_INV_RegFile[21][15]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux75~18_combout\,
	datag => \ALT_INV_RegFile[20][15]~q\,
	combout => \Mux75~5_combout\);

-- Location: MLABCELL_X72_Y2_N33
\Mux75~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux75~13_combout\ = ( \Mux75~26_combout\ & ( \Mux75~5_combout\ & ( (!\R.curInst\(18)) # ((!\R.curInst\(19) & ((\Mux75~1_combout\))) # (\R.curInst\(19) & (\Mux75~9_combout\))) ) ) ) # ( !\Mux75~26_combout\ & ( \Mux75~5_combout\ & ( (!\R.curInst\(19) & 
-- (\R.curInst\(18) & ((\Mux75~1_combout\)))) # (\R.curInst\(19) & ((!\R.curInst\(18)) # ((\Mux75~9_combout\)))) ) ) ) # ( \Mux75~26_combout\ & ( !\Mux75~5_combout\ & ( (!\R.curInst\(19) & ((!\R.curInst\(18)) # ((\Mux75~1_combout\)))) # (\R.curInst\(19) & 
-- (\R.curInst\(18) & (\Mux75~9_combout\))) ) ) ) # ( !\Mux75~26_combout\ & ( !\Mux75~5_combout\ & ( (\R.curInst\(18) & ((!\R.curInst\(19) & ((\Mux75~1_combout\))) # (\R.curInst\(19) & (\Mux75~9_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000100100011100010011010101101000101011001111100110111101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(19),
	datab => \ALT_INV_R.curInst\(18),
	datac => \ALT_INV_Mux75~9_combout\,
	datad => \ALT_INV_Mux75~1_combout\,
	datae => \ALT_INV_Mux75~26_combout\,
	dataf => \ALT_INV_Mux75~5_combout\,
	combout => \Mux75~13_combout\);

-- Location: LABCELL_X73_Y6_N54
\Mux239~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux239~0_combout\ = ( \Mux75~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC\(15)))) ) ) # ( !\Mux75~13_combout\ & ( (\R.curPC\(15) & (\vAluSrc1~2_combout\ & !\vAluSrc1~1_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000000000000110000000011110011000000001111001100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.curPC\(15),
	datac => \ALT_INV_vAluSrc1~2_combout\,
	datad => \ALT_INV_vAluSrc1~1_combout\,
	dataf => \ALT_INV_Mux75~13_combout\,
	combout => \Mux239~0_combout\);

-- Location: FF_X73_Y6_N16
\R.aluData1[15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux239~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData1\(15));

-- Location: LABCELL_X75_Y4_N27
\Mux140~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux140~0_combout\ = ( \Mux123~2_combout\ & ( \R.curInst\(14) ) ) # ( !\Mux123~2_combout\ & ( \R.curInst\(14) & ( ((\vAluSrc1~0_combout\ & ((\R.curInst\(2)) # (\Mux124~0_combout\)))) # (\Mux149~0_combout\) ) ) ) # ( \Mux123~2_combout\ & ( !\R.curInst\(14) 
-- ) ) # ( !\Mux123~2_combout\ & ( !\R.curInst\(14) & ( (\Mux124~0_combout\ & \vAluSrc1~0_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101111111111111111100000111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux124~0_combout\,
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_vAluSrc1~0_combout\,
	datad => \ALT_INV_Mux149~0_combout\,
	datae => \ALT_INV_Mux123~2_combout\,
	dataf => \ALT_INV_R.curInst\(14),
	combout => \Mux140~0_combout\);

-- Location: LABCELL_X80_Y3_N33
\R.regWriteData[14]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.regWriteData[14]~feeder_combout\ = \Add0~49_sumout\

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Add0~49_sumout\,
	combout => \R.regWriteData[14]~feeder_combout\);

-- Location: FF_X73_Y6_N34
\Add2~57_OTERM707_NEW_REG812\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux240~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Add2~57_OTERM707_OTERM813\);

-- Location: FF_X74_Y6_N4
\R.aluData1[13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux241~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData1\(13));

-- Location: LABCELL_X75_Y4_N51
\Mux142~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux142~0_combout\ = ( \Mux123~2_combout\ & ( \R.curInst\(12) ) ) # ( !\Mux123~2_combout\ & ( \R.curInst\(12) & ( ((\vAluSrc1~0_combout\ & ((\R.curInst\(2)) # (\Mux124~0_combout\)))) # (\Mux149~0_combout\) ) ) ) # ( \Mux123~2_combout\ & ( !\R.curInst\(12) 
-- ) ) # ( !\Mux123~2_combout\ & ( !\R.curInst\(12) & ( (\Mux124~0_combout\ & \vAluSrc1~0_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101111111111111111100000111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux124~0_combout\,
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_vAluSrc1~0_combout\,
	datad => \ALT_INV_Mux149~0_combout\,
	datae => \ALT_INV_Mux123~2_combout\,
	dataf => \ALT_INV_R.curInst\(12),
	combout => \Mux142~0_combout\);

-- Location: FF_X65_Y4_N2
\RegFile[31][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(12),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][12]~q\);

-- Location: FF_X68_Y6_N44
\RegFile[29][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(12),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][12]~q\);

-- Location: FF_X66_Y6_N43
\RegFile[30][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(12),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][12]~q\);

-- Location: FF_X65_Y4_N38
\RegFile[25][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(12),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][12]~q\);

-- Location: LABCELL_X57_Y4_N39
\RegFile[26][12]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[26][12]~feeder_combout\ = ( \R.regWriteData\(12) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(12),
	combout => \RegFile[26][12]~feeder_combout\);

-- Location: FF_X57_Y4_N40
\RegFile[26][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[26][12]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][12]~q\);

-- Location: FF_X65_Y4_N50
\RegFile[27][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(12),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][12]~q\);

-- Location: LABCELL_X57_Y4_N6
\RegFile[24][12]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[24][12]~feeder_combout\ = ( \R.regWriteData\(12) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(12),
	combout => \RegFile[24][12]~feeder_combout\);

-- Location: FF_X57_Y4_N7
\RegFile[24][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[24][12]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][12]~q\);

-- Location: MLABCELL_X65_Y4_N36
\Mux110~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux110~22_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[24][12]~q\))) # (\R.curInst\(20) & (\RegFile[25][12]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & (\RegFile[26][12]~q\)) # (\R.curInst\(20) & ((\RegFile[27][12]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[25][12]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[26][12]~q\,
	datad => \ALT_INV_RegFile[27][12]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][12]~q\,
	combout => \Mux110~22_combout\);

-- Location: MLABCELL_X65_Y9_N0
\RegFile[28][12]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[28][12]~feeder_combout\ = ( \R.regWriteData\(12) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(12),
	combout => \RegFile[28][12]~feeder_combout\);

-- Location: FF_X65_Y9_N1
\RegFile[28][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[28][12]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][12]~q\);

-- Location: LABCELL_X68_Y6_N42
\Mux110~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux110~9_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux110~22_combout\)))) # (\R.curInst\(22) & ((!\Mux110~22_combout\ & ((\RegFile[28][12]~q\))) # (\Mux110~22_combout\ & (\RegFile[29][12]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux110~22_combout\)))) # (\R.curInst\(22) & ((!\Mux110~22_combout\ & ((\RegFile[30][12]~q\))) # (\Mux110~22_combout\ & (\RegFile[31][12]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][12]~q\,
	datab => \ALT_INV_RegFile[29][12]~q\,
	datac => \ALT_INV_RegFile[30][12]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux110~22_combout\,
	datag => \ALT_INV_RegFile[28][12]~q\,
	combout => \Mux110~9_combout\);

-- Location: LABCELL_X64_Y9_N39
\RegFile[3][12]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[3][12]~feeder_combout\ = ( \R.regWriteData\(12) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(12),
	combout => \RegFile[3][12]~feeder_combout\);

-- Location: FF_X64_Y9_N40
\RegFile[3][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[3][12]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][12]~q\);

-- Location: FF_X65_Y6_N56
\RegFile[2][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(12),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][12]~q\);

-- Location: FF_X61_Y6_N41
\RegFile[5][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(12),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][12]~q\);

-- Location: FF_X65_Y6_N2
\RegFile[7][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(12),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][12]~q\);

-- Location: FF_X56_Y6_N8
\RegFile[4][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(12),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][12]~q\);

-- Location: FF_X65_Y6_N32
\RegFile[6][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(12),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][12]~q\);

-- Location: MLABCELL_X65_Y6_N30
\Mux110~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux110~0_combout\ = ( \RegFile[6][12]~q\ & ( \R.curInst\(21) & ( (!\R.curInst\(20)) # (\RegFile[7][12]~q\) ) ) ) # ( !\RegFile[6][12]~q\ & ( \R.curInst\(21) & ( (\RegFile[7][12]~q\ & \R.curInst\(20)) ) ) ) # ( \RegFile[6][12]~q\ & ( !\R.curInst\(21) & ( 
-- (!\R.curInst\(20) & ((\RegFile[4][12]~q\))) # (\R.curInst\(20) & (\RegFile[5][12]~q\)) ) ) ) # ( !\RegFile[6][12]~q\ & ( !\R.curInst\(21) & ( (!\R.curInst\(20) & ((\RegFile[4][12]~q\))) # (\R.curInst\(20) & (\RegFile[5][12]~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010111110101000001011111010100000011000000111111001111110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[5][12]~q\,
	datab => \ALT_INV_RegFile[7][12]~q\,
	datac => \ALT_INV_R.curInst\(20),
	datad => \ALT_INV_RegFile[4][12]~q\,
	datae => \ALT_INV_RegFile[6][12]~q\,
	dataf => \ALT_INV_R.curInst\(21),
	combout => \Mux110~0_combout\);

-- Location: LABCELL_X68_Y9_N57
\RegFile[1][12]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[1][12]~feeder_combout\ = ( \R.regWriteData\(12) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(12),
	combout => \RegFile[1][12]~feeder_combout\);

-- Location: FF_X68_Y9_N58
\RegFile[1][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[1][12]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][12]~q\);

-- Location: MLABCELL_X65_Y5_N36
\Mux110~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux110~26_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (\R.curInst\(20) & (\RegFile[1][12]~q\))) # (\R.curInst\(22) & (((\Mux110~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (((\RegFile[2][12]~q\)))) # 
-- (\R.curInst\(20) & (\RegFile[3][12]~q\)))) # (\R.curInst\(22) & ((((\Mux110~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000000000111010000000000000011111111110001110111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][12]~q\,
	datab => \ALT_INV_R.curInst\(20),
	datac => \ALT_INV_RegFile[2][12]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux110~0_combout\,
	datag => \ALT_INV_RegFile[1][12]~q\,
	combout => \Mux110~26_combout\);

-- Location: FF_X72_Y8_N52
\RegFile[21][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(12),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][12]~q\);

-- Location: FF_X70_Y8_N38
\RegFile[23][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(12),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][12]~q\);

-- Location: FF_X61_Y8_N58
\RegFile[22][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(12),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][12]~q\);

-- Location: FF_X64_Y8_N56
\RegFile[17][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(12),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][12]~q\);

-- Location: LABCELL_X71_Y4_N15
\RegFile[18][12]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[18][12]~feeder_combout\ = ( \R.regWriteData\(12) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(12),
	combout => \RegFile[18][12]~feeder_combout\);

-- Location: FF_X71_Y4_N16
\RegFile[18][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][12]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][12]~q\);

-- Location: FF_X70_Y4_N55
\RegFile[19][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(12),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][12]~q\);

-- Location: FF_X51_Y8_N25
\RegFile[16][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(12),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][12]~q\);

-- Location: LABCELL_X64_Y8_N54
\Mux110~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux110~18_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[16][12]~q\))) # (\R.curInst\(20) & (\RegFile[17][12]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & (\RegFile[18][12]~q\)) # (\R.curInst\(20) & ((\RegFile[19][12]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[17][12]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[18][12]~q\,
	datad => \ALT_INV_RegFile[19][12]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][12]~q\,
	combout => \Mux110~18_combout\);

-- Location: LABCELL_X60_Y8_N9
\RegFile[20][12]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[20][12]~feeder_combout\ = ( \R.regWriteData\(12) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(12),
	combout => \RegFile[20][12]~feeder_combout\);

-- Location: FF_X60_Y8_N10
\RegFile[20][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[20][12]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][12]~q\);

-- Location: LABCELL_X71_Y8_N12
\Mux110~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux110~5_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux110~18_combout\)))) # (\R.curInst\(22) & ((!\Mux110~18_combout\ & ((\RegFile[20][12]~q\))) # (\Mux110~18_combout\ & (\RegFile[21][12]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux110~18_combout\)))) # (\R.curInst\(22) & ((!\Mux110~18_combout\ & ((\RegFile[22][12]~q\))) # (\Mux110~18_combout\ & (\RegFile[23][12]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][12]~q\,
	datab => \ALT_INV_RegFile[23][12]~q\,
	datac => \ALT_INV_RegFile[22][12]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux110~18_combout\,
	datag => \ALT_INV_RegFile[20][12]~q\,
	combout => \Mux110~5_combout\);

-- Location: FF_X66_Y8_N44
\RegFile[15][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(12),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][12]~q\);

-- Location: FF_X61_Y8_N13
\RegFile[14][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(12),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][12]~q\);

-- Location: FF_X66_Y8_N26
\RegFile[9][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(12),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][12]~q\);

-- Location: LABCELL_X60_Y8_N21
\RegFile[10][12]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[10][12]~feeder_combout\ = ( \R.regWriteData\(12) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(12),
	combout => \RegFile[10][12]~feeder_combout\);

-- Location: FF_X60_Y8_N22
\RegFile[10][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[10][12]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][12]~q\);

-- Location: FF_X66_Y8_N8
\RegFile[11][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(12),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][12]~q\);

-- Location: FF_X63_Y8_N41
\RegFile[8][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(12),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][12]~q\);

-- Location: LABCELL_X66_Y8_N24
\Mux110~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux110~14_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[8][12]~q\))) # (\R.curInst\(20) & (\RegFile[9][12]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & (\RegFile[10][12]~q\)) # (\R.curInst\(20) & ((\RegFile[11][12]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][12]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[10][12]~q\,
	datad => \ALT_INV_RegFile[11][12]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][12]~q\,
	combout => \Mux110~14_combout\);

-- Location: LABCELL_X60_Y8_N24
\RegFile[12][12]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[12][12]~feeder_combout\ = ( \R.regWriteData\(12) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(12),
	combout => \RegFile[12][12]~feeder_combout\);

-- Location: FF_X60_Y8_N25
\RegFile[12][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[12][12]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][12]~q\);

-- Location: LABCELL_X66_Y8_N36
\Mux110~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux110~1_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux110~14_combout\)))) # (\R.curInst\(22) & ((!\Mux110~14_combout\ & ((\RegFile[12][12]~q\))) # (\Mux110~14_combout\ & (\RegFile[13][12]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux110~14_combout\)))) # (\R.curInst\(22) & ((!\Mux110~14_combout\ & ((\RegFile[14][12]~q\))) # (\Mux110~14_combout\ & (\RegFile[15][12]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][12]~q\,
	datab => \ALT_INV_RegFile[15][12]~q\,
	datac => \ALT_INV_RegFile[14][12]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux110~14_combout\,
	datag => \ALT_INV_RegFile[12][12]~q\,
	combout => \Mux110~1_combout\);

-- Location: LABCELL_X71_Y6_N48
\Mux110~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux110~13_combout\ = ( \Mux110~5_combout\ & ( \Mux110~1_combout\ & ( (!\R.curInst\(24) & (((\Mux110~26_combout\) # (\R.curInst\(23))))) # (\R.curInst\(24) & (((!\R.curInst\(23))) # (\Mux110~9_combout\))) ) ) ) # ( !\Mux110~5_combout\ & ( 
-- \Mux110~1_combout\ & ( (!\R.curInst\(24) & (((\Mux110~26_combout\) # (\R.curInst\(23))))) # (\R.curInst\(24) & (\Mux110~9_combout\ & (\R.curInst\(23)))) ) ) ) # ( \Mux110~5_combout\ & ( !\Mux110~1_combout\ & ( (!\R.curInst\(24) & (((!\R.curInst\(23) & 
-- \Mux110~26_combout\)))) # (\R.curInst\(24) & (((!\R.curInst\(23))) # (\Mux110~9_combout\))) ) ) ) # ( !\Mux110~5_combout\ & ( !\Mux110~1_combout\ & ( (!\R.curInst\(24) & (((!\R.curInst\(23) & \Mux110~26_combout\)))) # (\R.curInst\(24) & 
-- (\Mux110~9_combout\ & (\R.curInst\(23)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000111000001001100011111000100001101110011010011110111111101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux110~9_combout\,
	datab => \ALT_INV_R.curInst\(24),
	datac => \ALT_INV_R.curInst\(23),
	datad => \ALT_INV_Mux110~26_combout\,
	datae => \ALT_INV_Mux110~5_combout\,
	dataf => \ALT_INV_Mux110~1_combout\,
	combout => \Mux110~13_combout\);

-- Location: LABCELL_X71_Y6_N42
\NxR.aluData2[12]~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[12]~11_combout\ = ( \Mux110~13_combout\ & ( (!\vAluSrc2~1_combout\) # ((\Equal4~1_combout\ & \Mux142~0_combout\)) ) ) # ( !\Mux110~13_combout\ & ( (\Equal4~1_combout\ & (\vAluSrc2~1_combout\ & \Mux142~0_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000011000000000000001111110000111100111111000011110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Equal4~1_combout\,
	datac => \ALT_INV_vAluSrc2~1_combout\,
	datad => \ALT_INV_Mux142~0_combout\,
	dataf => \ALT_INV_Mux110~13_combout\,
	combout => \NxR.aluData2[12]~11_combout\);

-- Location: FF_X71_Y6_N58
\R.aluData2[12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \NxR.aluData2[12]~11_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData2\(12));

-- Location: LABCELL_X77_Y1_N18
\Mux143~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux143~0_combout\ = ( \R.curInst\(20) & ( (!\R.curInst\(2) & (\R.curInst\(7) & ((!\R.curInst\(3))))) # (\R.curInst\(2) & (((\R.curInst\(3)) # (\R.curInst\(31))))) ) ) # ( !\R.curInst\(20) & ( (!\R.curInst\(3) & ((!\R.curInst\(2) & (\R.curInst\(7))) # 
-- (\R.curInst\(2) & ((\R.curInst\(31)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101001100000000010100110000000001010011000011110101001100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(7),
	datab => \ALT_INV_R.curInst\(31),
	datac => \ALT_INV_R.curInst\(2),
	datad => \ALT_INV_R.curInst\(3),
	dataf => \ALT_INV_R.curInst\(20),
	combout => \Mux143~0_combout\);

-- Location: LABCELL_X77_Y1_N42
\Mux143~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux143~1_combout\ = ( \R.curInst\(4) & ( \Mux143~0_combout\ & ( (!\R.curInst\(6) & (\Mux53~0_combout\ & (!\R.curInst\(5) & \R.curInst\(31)))) ) ) ) # ( !\R.curInst\(4) & ( \Mux143~0_combout\ & ( (!\R.curInst\(6) & (\Mux53~0_combout\ & 
-- ((\R.curInst\(31))))) # (\R.curInst\(6) & (((\R.curInst\(5))))) ) ) ) # ( \R.curInst\(4) & ( !\Mux143~0_combout\ & ( (!\R.curInst\(6) & (\Mux53~0_combout\ & (!\R.curInst\(5) & \R.curInst\(31)))) ) ) ) # ( !\R.curInst\(4) & ( !\Mux143~0_combout\ & ( 
-- (!\R.curInst\(6) & (\Mux53~0_combout\ & \R.curInst\(31))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000100010000000000010000000000101001001110000000000100000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(6),
	datab => \ALT_INV_Mux53~0_combout\,
	datac => \ALT_INV_R.curInst\(5),
	datad => \ALT_INV_R.curInst\(31),
	datae => \ALT_INV_R.curInst\(4),
	dataf => \ALT_INV_Mux143~0_combout\,
	combout => \Mux143~1_combout\);

-- Location: FF_X73_Y2_N56
\RegFile[31][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(11),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][11]~q\);

-- Location: FF_X73_Y2_N13
\RegFile[30][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(11),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][11]~q\);

-- Location: FF_X67_Y2_N26
\RegFile[25][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(11),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][11]~q\);

-- Location: LABCELL_X67_Y2_N36
\RegFile[27][11]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[27][11]~feeder_combout\ = ( \R.regWriteData\(11) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(11),
	combout => \RegFile[27][11]~feeder_combout\);

-- Location: FF_X67_Y2_N37
\RegFile[27][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[27][11]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][11]~q\);

-- Location: LABCELL_X67_Y2_N33
\RegFile[26][11]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[26][11]~feeder_combout\ = ( \R.regWriteData\(11) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(11),
	combout => \RegFile[26][11]~feeder_combout\);

-- Location: FF_X67_Y2_N34
\RegFile[26][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[26][11]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][11]~q\);

-- Location: LABCELL_X56_Y2_N30
\RegFile[24][11]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[24][11]~feeder_combout\ = ( \R.regWriteData\(11) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(11),
	combout => \RegFile[24][11]~feeder_combout\);

-- Location: FF_X56_Y2_N31
\RegFile[24][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[24][11]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][11]~q\);

-- Location: LABCELL_X67_Y2_N24
\Mux111~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux111~22_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[24][11]~q\))) # (\R.curInst\(20) & (\RegFile[25][11]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[26][11]~q\))) # (\R.curInst\(20) & (\RegFile[27][11]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[25][11]~q\,
	datab => \ALT_INV_RegFile[27][11]~q\,
	datac => \ALT_INV_RegFile[26][11]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][11]~q\,
	combout => \Mux111~22_combout\);

-- Location: LABCELL_X73_Y2_N45
\RegFile[28][11]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[28][11]~feeder_combout\ = ( \R.regWriteData\(11) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(11),
	combout => \RegFile[28][11]~feeder_combout\);

-- Location: FF_X73_Y2_N47
\RegFile[28][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[28][11]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][11]~q\);

-- Location: LABCELL_X67_Y2_N12
\Mux111~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux111~9_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux111~22_combout\)))) # (\R.curInst\(22) & ((!\Mux111~22_combout\ & ((\RegFile[28][11]~q\))) # (\Mux111~22_combout\ & (\RegFile[29][11]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux111~22_combout\)))) # (\R.curInst\(22) & ((!\Mux111~22_combout\ & ((\RegFile[30][11]~q\))) # (\Mux111~22_combout\ & (\RegFile[31][11]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[29][11]~q\,
	datab => \ALT_INV_RegFile[31][11]~q\,
	datac => \ALT_INV_RegFile[30][11]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux111~22_combout\,
	datag => \ALT_INV_RegFile[28][11]~q\,
	combout => \Mux111~9_combout\);

-- Location: LABCELL_X70_Y2_N6
\RegFile[15][11]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[15][11]~feeder_combout\ = ( \R.regWriteData\(11) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(11),
	combout => \RegFile[15][11]~feeder_combout\);

-- Location: FF_X70_Y2_N7
\RegFile[15][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[15][11]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][11]~q\);

-- Location: FF_X74_Y2_N14
\RegFile[13][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(11),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][11]~q\);

-- Location: LABCELL_X62_Y2_N39
\RegFile[14][11]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[14][11]~feeder_combout\ = \R.regWriteData\(11)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.regWriteData\(11),
	combout => \RegFile[14][11]~feeder_combout\);

-- Location: FF_X62_Y2_N40
\RegFile[14][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[14][11]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][11]~q\);

-- Location: FF_X74_Y2_N50
\RegFile[9][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(11),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][11]~q\);

-- Location: LABCELL_X70_Y2_N42
\RegFile[11][11]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[11][11]~feeder_combout\ = ( \R.regWriteData\(11) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(11),
	combout => \RegFile[11][11]~feeder_combout\);

-- Location: FF_X70_Y2_N43
\RegFile[11][11]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[11][11]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][11]~DUPLICATE_q\);

-- Location: LABCELL_X75_Y2_N33
\RegFile[10][11]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[10][11]~feeder_combout\ = ( \R.regWriteData\(11) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(11),
	combout => \RegFile[10][11]~feeder_combout\);

-- Location: FF_X75_Y2_N34
\RegFile[10][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[10][11]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][11]~q\);

-- Location: LABCELL_X56_Y2_N3
\RegFile[8][11]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[8][11]~feeder_combout\ = ( \R.regWriteData\(11) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(11),
	combout => \RegFile[8][11]~feeder_combout\);

-- Location: FF_X56_Y2_N4
\RegFile[8][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[8][11]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][11]~q\);

-- Location: MLABCELL_X72_Y2_N48
\Mux111~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux111~14_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[8][11]~q\))) # (\R.curInst\(20) & (\RegFile[9][11]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[10][11]~q\))) # (\R.curInst\(20) & (\RegFile[11][11]~DUPLICATE_q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][11]~q\,
	datab => \ALT_INV_RegFile[11][11]~DUPLICATE_q\,
	datac => \ALT_INV_RegFile[10][11]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][11]~q\,
	combout => \Mux111~14_combout\);

-- Location: FF_X62_Y2_N28
\RegFile[12][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(11),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][11]~q\);

-- Location: LABCELL_X74_Y2_N12
\Mux111~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux111~1_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux111~14_combout\)))) # (\R.curInst\(22) & ((!\Mux111~14_combout\ & ((\RegFile[12][11]~q\))) # (\Mux111~14_combout\ & (\RegFile[13][11]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux111~14_combout\)))) # (\R.curInst\(22) & ((!\Mux111~14_combout\ & ((\RegFile[14][11]~q\))) # (\Mux111~14_combout\ & (\RegFile[15][11]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][11]~q\,
	datab => \ALT_INV_RegFile[13][11]~q\,
	datac => \ALT_INV_RegFile[14][11]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux111~14_combout\,
	datag => \ALT_INV_RegFile[12][11]~q\,
	combout => \Mux111~1_combout\);

-- Location: FF_X71_Y1_N2
\RegFile[21][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(11),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][11]~q\);

-- Location: FF_X72_Y1_N14
\RegFile[23][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(11),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][11]~q\);

-- Location: LABCELL_X71_Y1_N27
\RegFile[22][11]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[22][11]~feeder_combout\ = ( \R.regWriteData\(11) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(11),
	combout => \RegFile[22][11]~feeder_combout\);

-- Location: FF_X71_Y1_N29
\RegFile[22][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[22][11]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][11]~q\);

-- Location: FF_X72_Y1_N20
\RegFile[19][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(11),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][11]~q\);

-- Location: FF_X64_Y1_N38
\RegFile[17][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(11),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][11]~q\);

-- Location: FF_X73_Y1_N11
\RegFile[18][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(11),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][11]~q\);

-- Location: FF_X79_Y1_N5
\RegFile[16][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(11),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][11]~q\);

-- Location: LABCELL_X73_Y1_N9
\Mux111~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux111~18_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[16][11]~q\))) # (\R.curInst\(20) & (\RegFile[17][11]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[18][11]~q\))) # (\R.curInst\(20) & (\RegFile[19][11]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[19][11]~q\,
	datab => \ALT_INV_RegFile[17][11]~q\,
	datac => \ALT_INV_RegFile[18][11]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][11]~q\,
	combout => \Mux111~18_combout\);

-- Location: LABCELL_X75_Y1_N12
\RegFile[20][11]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[20][11]~feeder_combout\ = ( \R.regWriteData\(11) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(11),
	combout => \RegFile[20][11]~feeder_combout\);

-- Location: FF_X75_Y1_N13
\RegFile[20][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[20][11]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][11]~q\);

-- Location: LABCELL_X71_Y1_N0
\Mux111~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux111~5_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux111~18_combout\)))) # (\R.curInst\(22) & ((!\Mux111~18_combout\ & ((\RegFile[20][11]~q\))) # (\Mux111~18_combout\ & (\RegFile[21][11]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux111~18_combout\)))) # (\R.curInst\(22) & ((!\Mux111~18_combout\ & ((\RegFile[22][11]~q\))) # (\Mux111~18_combout\ & (\RegFile[23][11]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][11]~q\,
	datab => \ALT_INV_RegFile[23][11]~q\,
	datac => \ALT_INV_RegFile[22][11]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux111~18_combout\,
	datag => \ALT_INV_RegFile[20][11]~q\,
	combout => \Mux111~5_combout\);

-- Location: FF_X61_Y2_N20
\RegFile[3][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(11),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][11]~q\);

-- Location: FF_X62_Y1_N23
\RegFile[2][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(11),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][11]~q\);

-- Location: FF_X57_Y3_N13
\RegFile[6][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(11),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][11]~q\);

-- Location: FF_X61_Y2_N49
\RegFile[7][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(11),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][11]~q\);

-- Location: LABCELL_X56_Y2_N27
\RegFile[4][11]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[4][11]~feeder_combout\ = ( \R.regWriteData\(11) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(11),
	combout => \RegFile[4][11]~feeder_combout\);

-- Location: FF_X56_Y2_N28
\RegFile[4][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[4][11]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][11]~q\);

-- Location: FF_X61_Y2_N8
\RegFile[5][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(11),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][11]~q\);

-- Location: LABCELL_X61_Y2_N6
\Mux111~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux111~0_combout\ = ( \RegFile[5][11]~q\ & ( \R.curInst\(21) & ( (!\R.curInst\(20) & (\RegFile[6][11]~q\)) # (\R.curInst\(20) & ((\RegFile[7][11]~q\))) ) ) ) # ( !\RegFile[5][11]~q\ & ( \R.curInst\(21) & ( (!\R.curInst\(20) & (\RegFile[6][11]~q\)) # 
-- (\R.curInst\(20) & ((\RegFile[7][11]~q\))) ) ) ) # ( \RegFile[5][11]~q\ & ( !\R.curInst\(21) & ( (\RegFile[4][11]~q\) # (\R.curInst\(20)) ) ) ) # ( !\RegFile[5][11]~q\ & ( !\R.curInst\(21) & ( (!\R.curInst\(20) & \RegFile[4][11]~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011110000000011111111111101010011010100110101001101010011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[6][11]~q\,
	datab => \ALT_INV_RegFile[7][11]~q\,
	datac => \ALT_INV_R.curInst\(20),
	datad => \ALT_INV_RegFile[4][11]~q\,
	datae => \ALT_INV_RegFile[5][11]~q\,
	dataf => \ALT_INV_R.curInst\(21),
	combout => \Mux111~0_combout\);

-- Location: LABCELL_X53_Y3_N39
\RegFile[1][11]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[1][11]~feeder_combout\ = ( \R.regWriteData\(11) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(11),
	combout => \RegFile[1][11]~feeder_combout\);

-- Location: FF_X53_Y3_N40
\RegFile[1][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[1][11]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][11]~q\);

-- Location: LABCELL_X62_Y1_N21
\Mux111~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux111~26_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (\RegFile[1][11]~q\ & (\R.curInst\(20)))) # (\R.curInst\(22) & (((\Mux111~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (((\RegFile[2][11]~q\)))) # 
-- (\R.curInst\(20) & (\RegFile[3][11]~q\)))) # (\R.curInst\(22) & ((((\Mux111~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001100000011000100010000110011001111110011111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][11]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[2][11]~q\,
	datad => \ALT_INV_R.curInst\(20),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux111~0_combout\,
	datag => \ALT_INV_RegFile[1][11]~q\,
	combout => \Mux111~26_combout\);

-- Location: LABCELL_X74_Y2_N18
\Mux111~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux111~13_combout\ = ( \Mux111~5_combout\ & ( \Mux111~26_combout\ & ( (!\R.curInst\(23)) # ((!\R.curInst\(24) & ((\Mux111~1_combout\))) # (\R.curInst\(24) & (\Mux111~9_combout\))) ) ) ) # ( !\Mux111~5_combout\ & ( \Mux111~26_combout\ & ( 
-- (!\R.curInst\(23) & (((!\R.curInst\(24))))) # (\R.curInst\(23) & ((!\R.curInst\(24) & ((\Mux111~1_combout\))) # (\R.curInst\(24) & (\Mux111~9_combout\)))) ) ) ) # ( \Mux111~5_combout\ & ( !\Mux111~26_combout\ & ( (!\R.curInst\(23) & (((\R.curInst\(24))))) 
-- # (\R.curInst\(23) & ((!\R.curInst\(24) & ((\Mux111~1_combout\))) # (\R.curInst\(24) & (\Mux111~9_combout\)))) ) ) ) # ( !\Mux111~5_combout\ & ( !\Mux111~26_combout\ & ( (\R.curInst\(23) & ((!\R.curInst\(24) & ((\Mux111~1_combout\))) # (\R.curInst\(24) & 
-- (\Mux111~9_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000101010001000010110101101110100001111100011010101111111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(23),
	datab => \ALT_INV_Mux111~9_combout\,
	datac => \ALT_INV_R.curInst\(24),
	datad => \ALT_INV_Mux111~1_combout\,
	datae => \ALT_INV_Mux111~5_combout\,
	dataf => \ALT_INV_Mux111~26_combout\,
	combout => \Mux111~13_combout\);

-- Location: LABCELL_X75_Y6_N12
\NxR.aluData2[11]~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[11]~8_combout\ = ( \Mux111~13_combout\ & ( (!\vAluSrc2~1_combout\) # ((\Equal4~1_combout\ & \Mux143~1_combout\)) ) ) # ( !\Mux111~13_combout\ & ( (\Equal4~1_combout\ & (\Mux143~1_combout\ & \vAluSrc2~1_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000101000000000000010111111111000001011111111100000101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Equal4~1_combout\,
	datac => \ALT_INV_Mux143~1_combout\,
	datad => \ALT_INV_vAluSrc2~1_combout\,
	dataf => \ALT_INV_Mux111~13_combout\,
	combout => \NxR.aluData2[11]~8_combout\);

-- Location: FF_X75_Y6_N44
\R.aluData2[11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \NxR.aluData2[11]~8_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData2\(11));

-- Location: FF_X75_Y6_N8
\Add2~41_OTERM715_NEW_REG818\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \NxR.aluData2[10]~9_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Add2~41_OTERM715_OTERM819\);

-- Location: LABCELL_X67_Y8_N18
\RegFile[13][10]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[13][10]~feeder_combout\ = ( \R.regWriteData\(10) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(10),
	combout => \RegFile[13][10]~feeder_combout\);

-- Location: FF_X67_Y8_N20
\RegFile[13][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[13][10]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][10]~q\);

-- Location: LABCELL_X67_Y8_N48
\RegFile[14][10]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[14][10]~feeder_combout\ = ( \R.regWriteData\(10) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(10),
	combout => \RegFile[14][10]~feeder_combout\);

-- Location: FF_X67_Y8_N49
\RegFile[14][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[14][10]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][10]~q\);

-- Location: FF_X66_Y7_N58
\RegFile[15][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(10),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][10]~q\);

-- Location: LABCELL_X68_Y8_N0
\RegFile[9][10]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[9][10]~feeder_combout\ = ( \R.regWriteData\(10) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(10),
	combout => \RegFile[9][10]~feeder_combout\);

-- Location: FF_X68_Y8_N1
\RegFile[9][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[9][10]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][10]~q\);

-- Location: FF_X64_Y8_N29
\RegFile[11][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(10),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][10]~q\);

-- Location: LABCELL_X60_Y8_N36
\RegFile[10][10]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[10][10]~feeder_combout\ = ( \R.regWriteData\(10) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(10),
	combout => \RegFile[10][10]~feeder_combout\);

-- Location: FF_X60_Y8_N38
\RegFile[10][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[10][10]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][10]~q\);

-- Location: LABCELL_X63_Y8_N3
\RegFile[8][10]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[8][10]~feeder_combout\ = ( \R.regWriteData\(10) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(10),
	combout => \RegFile[8][10]~feeder_combout\);

-- Location: FF_X63_Y8_N4
\RegFile[8][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[8][10]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][10]~q\);

-- Location: LABCELL_X64_Y8_N27
\Mux80~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux80~14_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[8][10]~q\))) # (\R.curInst\(15) & (\RegFile[9][10]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[10][10]~q\))) # (\R.curInst\(15) & (\RegFile[11][10]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][10]~q\,
	datab => \ALT_INV_RegFile[11][10]~q\,
	datac => \ALT_INV_RegFile[10][10]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][10]~q\,
	combout => \Mux80~14_combout\);

-- Location: LABCELL_X70_Y8_N0
\RegFile[12][10]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[12][10]~feeder_combout\ = ( \R.regWriteData\(10) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(10),
	combout => \RegFile[12][10]~feeder_combout\);

-- Location: FF_X70_Y8_N2
\RegFile[12][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[12][10]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][10]~q\);

-- Location: LABCELL_X73_Y8_N27
\Mux80~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux80~1_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux80~14_combout\))))) # (\R.curInst\(17) & (((!\Mux80~14_combout\ & ((\RegFile[12][10]~q\))) # (\Mux80~14_combout\ & (\RegFile[13][10]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux80~14_combout\)))) # (\R.curInst\(17) & ((!\Mux80~14_combout\ & (\RegFile[14][10]~q\)) # (\Mux80~14_combout\ & ((\RegFile[15][10]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][10]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[14][10]~q\,
	datad => \ALT_INV_RegFile[15][10]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux80~14_combout\,
	datag => \ALT_INV_RegFile[12][10]~q\,
	combout => \Mux80~1_combout\);

-- Location: FF_X64_Y6_N50
\RegFile[31][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(10),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][10]~q\);

-- Location: FF_X66_Y6_N26
\RegFile[30][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(10),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][10]~q\);

-- Location: FF_X66_Y6_N56
\RegFile[29][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(10),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][10]~q\);

-- Location: FF_X64_Y6_N32
\RegFile[27][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(10),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][10]~q\);

-- Location: FF_X60_Y6_N7
\RegFile[26][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(10),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][10]~q\);

-- Location: FF_X66_Y6_N14
\RegFile[25][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(10),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][10]~q\);

-- Location: FF_X64_Y6_N59
\RegFile[24][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(10),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][10]~q\);

-- Location: LABCELL_X64_Y6_N30
\Mux80~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux80~22_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & (\RegFile[24][10]~q\)) # (\R.curInst\(15) & ((\RegFile[25][10]~q\)))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & ((\RegFile[26][10]~q\))) # (\R.curInst\(15) & (\RegFile[27][10]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001010101111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[27][10]~q\,
	datac => \ALT_INV_RegFile[26][10]~q\,
	datad => \ALT_INV_RegFile[25][10]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][10]~q\,
	combout => \Mux80~22_combout\);

-- Location: FF_X60_Y6_N13
\RegFile[28][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(10),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][10]~q\);

-- Location: LABCELL_X64_Y6_N48
\Mux80~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux80~9_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux80~22_combout\))))) # (\R.curInst\(17) & (((!\Mux80~22_combout\ & (\RegFile[28][10]~q\)) # (\Mux80~22_combout\ & ((\RegFile[29][10]~q\)))))) ) ) # ( \R.curInst\(16) & ( 
-- (!\R.curInst\(17) & ((((\Mux80~22_combout\))))) # (\R.curInst\(17) & (((!\Mux80~22_combout\ & ((\RegFile[30][10]~q\))) # (\Mux80~22_combout\ & (\RegFile[31][10]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110101010111111111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[31][10]~q\,
	datac => \ALT_INV_RegFile[30][10]~q\,
	datad => \ALT_INV_RegFile[29][10]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux80~22_combout\,
	datag => \ALT_INV_RegFile[28][10]~q\,
	combout => \Mux80~9_combout\);

-- Location: FF_X65_Y8_N32
\RegFile[21][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(10),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][10]~q\);

-- Location: FF_X75_Y8_N13
\RegFile[23][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(10),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][10]~q\);

-- Location: FF_X75_Y8_N37
\RegFile[22][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(10),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][10]~q\);

-- Location: FF_X65_Y8_N26
\RegFile[17][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(10),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][10]~q\);

-- Location: FF_X64_Y10_N4
\RegFile[18][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(10),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][10]~q\);

-- Location: MLABCELL_X65_Y8_N12
\RegFile[19][10]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[19][10]~feeder_combout\ = ( \R.regWriteData\(10) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(10),
	combout => \RegFile[19][10]~feeder_combout\);

-- Location: FF_X65_Y8_N13
\RegFile[19][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[19][10]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][10]~q\);

-- Location: LABCELL_X63_Y9_N51
\RegFile[16][10]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[16][10]~feeder_combout\ = ( \R.regWriteData\(10) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(10),
	combout => \RegFile[16][10]~feeder_combout\);

-- Location: FF_X63_Y9_N52
\RegFile[16][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[16][10]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][10]~q\);

-- Location: LABCELL_X74_Y8_N6
\Mux80~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux80~18_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[16][10]~q\))) # (\R.curInst\(15) & (\RegFile[17][10]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & (\RegFile[18][10]~q\)) # (\R.curInst\(15) & ((\RegFile[19][10]~q\)))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001110111011101110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[17][10]~q\,
	datac => \ALT_INV_RegFile[18][10]~q\,
	datad => \ALT_INV_RegFile[19][10]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][10]~q\,
	combout => \Mux80~18_combout\);

-- Location: FF_X64_Y10_N40
\RegFile[20][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(10),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][10]~q\);

-- Location: LABCELL_X74_Y8_N36
\Mux80~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux80~5_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux80~18_combout\)))) # (\R.curInst\(17) & ((!\Mux80~18_combout\ & ((\RegFile[20][10]~q\))) # (\Mux80~18_combout\ & (\RegFile[21][10]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux80~18_combout\)))) # (\R.curInst\(17) & ((!\Mux80~18_combout\ & ((\RegFile[22][10]~q\))) # (\Mux80~18_combout\ & (\RegFile[23][10]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][10]~q\,
	datab => \ALT_INV_RegFile[23][10]~q\,
	datac => \ALT_INV_RegFile[22][10]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux80~18_combout\,
	datag => \ALT_INV_RegFile[20][10]~q\,
	combout => \Mux80~5_combout\);

-- Location: FF_X62_Y8_N38
\RegFile[3][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(10),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][10]~q\);

-- Location: FF_X65_Y6_N26
\RegFile[6][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(10),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][10]~q\);

-- Location: LABCELL_X62_Y8_N42
\RegFile[5][10]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[5][10]~feeder_combout\ = ( \R.regWriteData\(10) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(10),
	combout => \RegFile[5][10]~feeder_combout\);

-- Location: FF_X62_Y8_N43
\RegFile[5][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[5][10]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][10]~q\);

-- Location: FF_X62_Y8_N25
\RegFile[7][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(10),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][10]~q\);

-- Location: FF_X56_Y6_N37
\RegFile[4][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(10),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][10]~q\);

-- Location: LABCELL_X62_Y8_N24
\Mux80~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux80~0_combout\ = ( \RegFile[7][10]~q\ & ( \RegFile[4][10]~q\ & ( (!\R.curInst\(16) & (((!\R.curInst\(15)) # (\RegFile[5][10]~q\)))) # (\R.curInst\(16) & (((\R.curInst\(15))) # (\RegFile[6][10]~q\))) ) ) ) # ( !\RegFile[7][10]~q\ & ( \RegFile[4][10]~q\ 
-- & ( (!\R.curInst\(16) & (((!\R.curInst\(15)) # (\RegFile[5][10]~q\)))) # (\R.curInst\(16) & (\RegFile[6][10]~q\ & ((!\R.curInst\(15))))) ) ) ) # ( \RegFile[7][10]~q\ & ( !\RegFile[4][10]~q\ & ( (!\R.curInst\(16) & (((\RegFile[5][10]~q\ & 
-- \R.curInst\(15))))) # (\R.curInst\(16) & (((\R.curInst\(15))) # (\RegFile[6][10]~q\))) ) ) ) # ( !\RegFile[7][10]~q\ & ( !\RegFile[4][10]~q\ & ( (!\R.curInst\(16) & (((\RegFile[5][10]~q\ & \R.curInst\(15))))) # (\R.curInst\(16) & (\RegFile[6][10]~q\ & 
-- ((!\R.curInst\(15))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100110000000001010011111111110101001100001111010100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[6][10]~q\,
	datab => \ALT_INV_RegFile[5][10]~q\,
	datac => \ALT_INV_R.curInst\(16),
	datad => \ALT_INV_R.curInst\(15),
	datae => \ALT_INV_RegFile[7][10]~q\,
	dataf => \ALT_INV_RegFile[4][10]~q\,
	combout => \Mux80~0_combout\);

-- Location: MLABCELL_X59_Y7_N9
\RegFile[1][10]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[1][10]~feeder_combout\ = ( \R.regWriteData\(10) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(10),
	combout => \RegFile[1][10]~feeder_combout\);

-- Location: FF_X59_Y7_N10
\RegFile[1][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[1][10]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][10]~q\);

-- Location: LABCELL_X62_Y8_N36
\Mux80~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux80~26_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (\R.curInst\(15) & (\RegFile[1][10]~q\))) # (\R.curInst\(17) & (((\Mux80~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & ((!\R.curInst\(15) & (((\RegFile[2][10]~q\)))) # 
-- (\R.curInst\(15) & (\RegFile[3][10]~q\)))) # (\R.curInst\(17) & ((((\Mux80~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000000000111010000000000000011111111110001110111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][10]~q\,
	datab => \ALT_INV_R.curInst\(15),
	datac => \ALT_INV_RegFile[2][10]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux80~0_combout\,
	datag => \ALT_INV_RegFile[1][10]~q\,
	combout => \Mux80~26_combout\);

-- Location: LABCELL_X74_Y8_N30
\Mux80~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux80~13_combout\ = ( \Mux80~5_combout\ & ( \Mux80~26_combout\ & ( (!\R.curInst\(18)) # ((!\R.curInst\(19) & (\Mux80~1_combout\)) # (\R.curInst\(19) & ((\Mux80~9_combout\)))) ) ) ) # ( !\Mux80~5_combout\ & ( \Mux80~26_combout\ & ( (!\R.curInst\(19) & 
-- ((!\R.curInst\(18)) # ((\Mux80~1_combout\)))) # (\R.curInst\(19) & (\R.curInst\(18) & ((\Mux80~9_combout\)))) ) ) ) # ( \Mux80~5_combout\ & ( !\Mux80~26_combout\ & ( (!\R.curInst\(19) & (\R.curInst\(18) & (\Mux80~1_combout\))) # (\R.curInst\(19) & 
-- ((!\R.curInst\(18)) # ((\Mux80~9_combout\)))) ) ) ) # ( !\Mux80~5_combout\ & ( !\Mux80~26_combout\ & ( (\R.curInst\(18) & ((!\R.curInst\(19) & (\Mux80~1_combout\)) # (\R.curInst\(19) & ((\Mux80~9_combout\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001000010011010001100101011110001010100110111100111011011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(19),
	datab => \ALT_INV_R.curInst\(18),
	datac => \ALT_INV_Mux80~1_combout\,
	datad => \ALT_INV_Mux80~9_combout\,
	datae => \ALT_INV_Mux80~5_combout\,
	dataf => \ALT_INV_Mux80~26_combout\,
	combout => \Mux80~13_combout\);

-- Location: LABCELL_X74_Y8_N0
\Mux244~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux244~0_combout\ = ( \Mux80~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC\(10)))) ) ) # ( !\Mux80~13_combout\ & ( (\vAluSrc1~2_combout\ & (\R.curPC\(10) & !\vAluSrc1~1_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000000000000110000000011001111000000001100111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_vAluSrc1~2_combout\,
	datac => \ALT_INV_R.curPC\(10),
	datad => \ALT_INV_vAluSrc1~1_combout\,
	dataf => \ALT_INV_Mux80~13_combout\,
	combout => \Mux244~0_combout\);

-- Location: LABCELL_X75_Y8_N9
\Add2~41_OTERM715_OTERM817feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~41_OTERM715_OTERM817feeder_combout\ = ( \Mux244~0_combout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_Mux244~0_combout\,
	combout => \Add2~41_OTERM715_OTERM817feeder_combout\);

-- Location: FF_X75_Y8_N10
\Add2~41_OTERM715_NEW_REG816\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Add2~41_OTERM715_OTERM817feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Add2~41_OTERM715_OTERM817\);

-- Location: LABCELL_X77_Y1_N48
\Mux145~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux145~0_combout\ = ( \R.curInst\(29) & ( \R.curInst\(5) & ( (!\R.curInst\(4) & ((!\R.curInst\(2) & ((!\R.curInst\(3)))) # (\R.curInst\(2) & (\R.curInst\(6))))) ) ) ) # ( \R.curInst\(29) & ( !\R.curInst\(5) & ( (!\R.curInst\(2) & (!\R.curInst\(6) & 
-- !\R.curInst\(3))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101000000000000000000000000000001000110000000100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(2),
	datab => \ALT_INV_R.curInst\(4),
	datac => \ALT_INV_R.curInst\(6),
	datad => \ALT_INV_R.curInst\(3),
	datae => \ALT_INV_R.curInst\(29),
	dataf => \ALT_INV_R.curInst\(5),
	combout => \Mux145~0_combout\);

-- Location: LABCELL_X81_Y6_N18
\Add0~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~25_sumout\ = SUM(( \R.curPC\(8) ) + ( GND ) + ( \Add0~22\ ))
-- \Add0~26\ = CARRY(( \R.curPC\(8) ) + ( GND ) + ( \Add0~22\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \ALT_INV_R.curPC\(8),
	cin => \Add0~22\,
	sumout => \Add0~25_sumout\,
	cout => \Add0~26\);

-- Location: LABCELL_X81_Y6_N21
\Add0~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~29_sumout\ = SUM(( \R.curPC\(9) ) + ( GND ) + ( \Add0~26\ ))
-- \Add0~30\ = CARRY(( \R.curPC\(9) ) + ( GND ) + ( \Add0~26\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.curPC\(9),
	cin => \Add0~26\,
	sumout => \Add0~29_sumout\,
	cout => \Add0~30\);

-- Location: LABCELL_X80_Y3_N3
\R.regWriteData[9]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.regWriteData[9]~feeder_combout\ = ( \Add0~29_sumout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_Add0~29_sumout\,
	combout => \R.regWriteData[9]~feeder_combout\);

-- Location: LABCELL_X66_Y3_N48
\RegFile[31][9]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[31][9]~feeder_combout\ = ( \R.regWriteData\(9) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(9),
	combout => \RegFile[31][9]~feeder_combout\);

-- Location: FF_X66_Y3_N49
\RegFile[31][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[31][9]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][9]~q\);

-- Location: LABCELL_X66_Y3_N39
\RegFile[30][9]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[30][9]~feeder_combout\ = ( \R.regWriteData\(9) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(9),
	combout => \RegFile[30][9]~feeder_combout\);

-- Location: FF_X66_Y3_N40
\RegFile[30][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[30][9]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][9]~q\);

-- Location: LABCELL_X68_Y1_N30
\RegFile[29][9]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[29][9]~feeder_combout\ = ( \R.regWriteData\(9) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(9),
	combout => \RegFile[29][9]~feeder_combout\);

-- Location: FF_X68_Y1_N31
\RegFile[29][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[29][9]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][9]~q\);

-- Location: FF_X67_Y1_N14
\RegFile[25][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(9),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][9]~q\);

-- Location: LABCELL_X67_Y2_N30
\RegFile[26][9]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[26][9]~feeder_combout\ = \R.regWriteData\(9)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.regWriteData\(9),
	combout => \RegFile[26][9]~feeder_combout\);

-- Location: FF_X67_Y2_N31
\RegFile[26][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[26][9]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][9]~q\);

-- Location: FF_X64_Y6_N25
\RegFile[27][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(9),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][9]~q\);

-- Location: FF_X64_Y6_N43
\RegFile[24][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(9),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][9]~q\);

-- Location: LABCELL_X64_Y6_N0
\Mux81~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux81~22_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[24][9]~q\))) # (\R.curInst\(15) & (\RegFile[25][9]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & (\RegFile[26][9]~q\)) # (\R.curInst\(15) & ((\RegFile[27][9]~q\)))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001110111011101110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[25][9]~q\,
	datac => \ALT_INV_RegFile[26][9]~q\,
	datad => \ALT_INV_RegFile[27][9]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][9]~q\,
	combout => \Mux81~22_combout\);

-- Location: FF_X66_Y3_N22
\RegFile[28][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(9),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][9]~q\);

-- Location: MLABCELL_X65_Y6_N42
\Mux81~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux81~9_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux81~22_combout\)))) # (\R.curInst\(17) & ((!\Mux81~22_combout\ & (\RegFile[28][9]~q\)) # (\Mux81~22_combout\ & ((\RegFile[29][9]~q\)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- ((((\Mux81~22_combout\))))) # (\R.curInst\(17) & (((!\Mux81~22_combout\ & ((\RegFile[30][9]~q\))) # (\Mux81~22_combout\ & (\RegFile[31][9]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111001100111111111101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][9]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[30][9]~q\,
	datad => \ALT_INV_RegFile[29][9]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux81~22_combout\,
	datag => \ALT_INV_RegFile[28][9]~q\,
	combout => \Mux81~9_combout\);

-- Location: FF_X65_Y5_N19
\RegFile[14][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(9),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][9]~q\);

-- Location: FF_X65_Y5_N38
\RegFile[15][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(9),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][9]~q\);

-- Location: FF_X64_Y3_N14
\RegFile[9][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(9),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][9]~q\);

-- Location: FF_X64_Y3_N23
\RegFile[10][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(9),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][9]~q\);

-- Location: FF_X64_Y3_N44
\RegFile[11][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(9),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][9]~q\);

-- Location: LABCELL_X66_Y5_N36
\RegFile[8][9]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[8][9]~feeder_combout\ = ( \R.regWriteData\(9) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(9),
	combout => \RegFile[8][9]~feeder_combout\);

-- Location: FF_X66_Y5_N37
\RegFile[8][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[8][9]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][9]~q\);

-- Location: LABCELL_X64_Y3_N42
\Mux81~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux81~14_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[8][9]~q\))) # (\R.curInst\(15) & (\RegFile[9][9]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & (\RegFile[10][9]~q\)) # (\R.curInst\(15) & ((\RegFile[11][9]~q\)))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001110111011101110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[9][9]~q\,
	datac => \ALT_INV_RegFile[10][9]~q\,
	datad => \ALT_INV_RegFile[11][9]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][9]~q\,
	combout => \Mux81~14_combout\);

-- Location: LABCELL_X60_Y5_N30
\RegFile[12][9]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[12][9]~feeder_combout\ = ( \R.regWriteData\(9) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(9),
	combout => \RegFile[12][9]~feeder_combout\);

-- Location: FF_X60_Y5_N31
\RegFile[12][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[12][9]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][9]~q\);

-- Location: MLABCELL_X65_Y6_N36
\Mux81~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux81~1_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux81~14_combout\))))) # (\R.curInst\(17) & (((!\Mux81~14_combout\ & ((\RegFile[12][9]~q\))) # (\Mux81~14_combout\ & (\RegFile[13][9]~q\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) 
-- & ((((\Mux81~14_combout\))))) # (\R.curInst\(17) & (((!\Mux81~14_combout\ & (\RegFile[14][9]~q\)) # (\Mux81~14_combout\ & ((\RegFile[15][9]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110111011101110111010101011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[13][9]~q\,
	datac => \ALT_INV_RegFile[14][9]~q\,
	datad => \ALT_INV_RegFile[15][9]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux81~14_combout\,
	datag => \ALT_INV_RegFile[12][9]~q\,
	combout => \Mux81~1_combout\);

-- Location: FF_X64_Y4_N20
\RegFile[23][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(9),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][9]~q\);

-- Location: FF_X64_Y5_N5
\RegFile[21][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(9),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][9]~q\);

-- Location: LABCELL_X64_Y4_N0
\RegFile[22][9]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[22][9]~feeder_combout\ = \R.regWriteData\(9)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.regWriteData\(9),
	combout => \RegFile[22][9]~feeder_combout\);

-- Location: FF_X64_Y4_N2
\RegFile[22][9]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[22][9]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][9]~DUPLICATE_q\);

-- Location: FF_X57_Y5_N10
\RegFile[17][9]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(9),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][9]~DUPLICATE_q\);

-- Location: LABCELL_X63_Y5_N9
\RegFile[18][9]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[18][9]~feeder_combout\ = ( \R.regWriteData\(9) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(9),
	combout => \RegFile[18][9]~feeder_combout\);

-- Location: FF_X63_Y5_N11
\RegFile[18][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][9]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][9]~q\);

-- Location: FF_X64_Y4_N8
\RegFile[19][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(9),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][9]~q\);

-- Location: LABCELL_X63_Y5_N39
\RegFile[16][9]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[16][9]~feeder_combout\ = \R.regWriteData\(9)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101010101010101010101010101010101010101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.regWriteData\(9),
	combout => \RegFile[16][9]~feeder_combout\);

-- Location: FF_X63_Y5_N41
\RegFile[16][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[16][9]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][9]~q\);

-- Location: LABCELL_X64_Y4_N6
\Mux81~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux81~18_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[16][9]~q\))) # (\R.curInst\(15) & (\RegFile[17][9]~DUPLICATE_q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( 
-- (!\R.curInst\(17) & (((!\R.curInst\(15) & (\RegFile[18][9]~q\)) # (\R.curInst\(15) & ((\RegFile[19][9]~q\)))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001110111011101110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[17][9]~DUPLICATE_q\,
	datac => \ALT_INV_RegFile[18][9]~q\,
	datad => \ALT_INV_RegFile[19][9]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][9]~q\,
	combout => \Mux81~18_combout\);

-- Location: FF_X59_Y4_N4
\RegFile[20][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(9),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][9]~q\);

-- Location: LABCELL_X64_Y4_N18
\Mux81~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux81~5_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux81~18_combout\)))) # (\R.curInst\(17) & ((!\Mux81~18_combout\ & ((\RegFile[20][9]~q\))) # (\Mux81~18_combout\ & (\RegFile[21][9]~q\))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) 
-- & (((\Mux81~18_combout\)))) # (\R.curInst\(17) & ((!\Mux81~18_combout\ & ((\RegFile[22][9]~DUPLICATE_q\))) # (\Mux81~18_combout\ & (\RegFile[23][9]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[23][9]~q\,
	datab => \ALT_INV_RegFile[21][9]~q\,
	datac => \ALT_INV_RegFile[22][9]~DUPLICATE_q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux81~18_combout\,
	datag => \ALT_INV_RegFile[20][9]~q\,
	combout => \Mux81~5_combout\);

-- Location: FF_X61_Y2_N38
\RegFile[3][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(9),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][9]~q\);

-- Location: FF_X61_Y5_N56
\RegFile[2][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(9),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][9]~q\);

-- Location: FF_X56_Y4_N19
\RegFile[6][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(9),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][9]~q\);

-- Location: FF_X61_Y2_N44
\RegFile[5][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(9),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][9]~q\);

-- Location: FF_X56_Y4_N13
\RegFile[4][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(9),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][9]~q\);

-- Location: FF_X61_Y2_N13
\RegFile[7][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(9),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][9]~q\);

-- Location: LABCELL_X61_Y2_N12
\Mux81~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux81~0_combout\ = ( \RegFile[7][9]~q\ & ( \R.curInst\(15) & ( (\R.curInst\(16)) # (\RegFile[5][9]~q\) ) ) ) # ( !\RegFile[7][9]~q\ & ( \R.curInst\(15) & ( (\RegFile[5][9]~q\ & !\R.curInst\(16)) ) ) ) # ( \RegFile[7][9]~q\ & ( !\R.curInst\(15) & ( 
-- (!\R.curInst\(16) & ((\RegFile[4][9]~q\))) # (\R.curInst\(16) & (\RegFile[6][9]~q\)) ) ) ) # ( !\RegFile[7][9]~q\ & ( !\R.curInst\(15) & ( (!\R.curInst\(16) & ((\RegFile[4][9]~q\))) # (\R.curInst\(16) & (\RegFile[6][9]~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010111110101000001011111010100110000001100000011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[6][9]~q\,
	datab => \ALT_INV_RegFile[5][9]~q\,
	datac => \ALT_INV_R.curInst\(16),
	datad => \ALT_INV_RegFile[4][9]~q\,
	datae => \ALT_INV_RegFile[7][9]~q\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux81~0_combout\);

-- Location: FF_X61_Y5_N44
\RegFile[1][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(9),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][9]~q\);

-- Location: LABCELL_X61_Y2_N36
\Mux81~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux81~26_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (\RegFile[1][9]~q\ & (\R.curInst\(15)))) # (\R.curInst\(17) & (((\Mux81~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & ((!\R.curInst\(15) & (((\RegFile[2][9]~q\)))) # 
-- (\R.curInst\(15) & (\RegFile[3][9]~q\)))) # (\R.curInst\(17) & ((((\Mux81~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001100000011000100010000110011001111110011111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][9]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[2][9]~q\,
	datad => \ALT_INV_R.curInst\(15),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux81~0_combout\,
	datag => \ALT_INV_RegFile[1][9]~q\,
	combout => \Mux81~26_combout\);

-- Location: MLABCELL_X65_Y6_N57
\Mux81~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux81~13_combout\ = ( \Mux81~5_combout\ & ( \Mux81~26_combout\ & ( (!\R.curInst\(18)) # ((!\R.curInst\(19) & ((\Mux81~1_combout\))) # (\R.curInst\(19) & (\Mux81~9_combout\))) ) ) ) # ( !\Mux81~5_combout\ & ( \Mux81~26_combout\ & ( (!\R.curInst\(19) & 
-- ((!\R.curInst\(18)) # ((\Mux81~1_combout\)))) # (\R.curInst\(19) & (\R.curInst\(18) & (\Mux81~9_combout\))) ) ) ) # ( \Mux81~5_combout\ & ( !\Mux81~26_combout\ & ( (!\R.curInst\(19) & (\R.curInst\(18) & ((\Mux81~1_combout\)))) # (\R.curInst\(19) & 
-- ((!\R.curInst\(18)) # ((\Mux81~9_combout\)))) ) ) ) # ( !\Mux81~5_combout\ & ( !\Mux81~26_combout\ & ( (\R.curInst\(18) & ((!\R.curInst\(19) & ((\Mux81~1_combout\))) # (\R.curInst\(19) & (\Mux81~9_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000100100011010001010110011110001001101010111100110111101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(19),
	datab => \ALT_INV_R.curInst\(18),
	datac => \ALT_INV_Mux81~9_combout\,
	datad => \ALT_INV_Mux81~1_combout\,
	datae => \ALT_INV_Mux81~5_combout\,
	dataf => \ALT_INV_Mux81~26_combout\,
	combout => \Mux81~13_combout\);

-- Location: LABCELL_X74_Y7_N57
\Mux245~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux245~0_combout\ = ( \Mux81~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC\(9)))) ) ) # ( !\Mux81~13_combout\ & ( (!\vAluSrc1~1_combout\ & (\vAluSrc1~2_combout\ & \R.curPC\(9))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001000000010000000100000001010001010100010101000101010001010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluSrc1~1_combout\,
	datab => \ALT_INV_vAluSrc1~2_combout\,
	datac => \ALT_INV_R.curPC\(9),
	dataf => \ALT_INV_Mux81~13_combout\,
	combout => \Mux245~0_combout\);

-- Location: FF_X78_Y7_N10
\Add2~33_OTERM719_NEW_REG820\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux245~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Add2~33_OTERM719_OTERM821\);

-- Location: FF_X62_Y6_N2
\RegFile[29][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(7),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][7]~q\);

-- Location: FF_X62_Y4_N2
\RegFile[31][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(7),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][7]~q\);

-- Location: LABCELL_X62_Y6_N6
\RegFile[30][7]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[30][7]~feeder_combout\ = ( \R.regWriteData\(7) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(7),
	combout => \RegFile[30][7]~feeder_combout\);

-- Location: FF_X62_Y6_N8
\RegFile[30][7]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[30][7]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][7]~DUPLICATE_q\);

-- Location: FF_X62_Y4_N32
\RegFile[25][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(7),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][7]~q\);

-- Location: FF_X57_Y3_N19
\RegFile[26][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(7),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][7]~q\);

-- Location: FF_X62_Y4_N26
\RegFile[27][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(7),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][7]~q\);

-- Location: LABCELL_X60_Y3_N48
\RegFile[24][7]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[24][7]~feeder_combout\ = ( \R.regWriteData\(7) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(7),
	combout => \RegFile[24][7]~feeder_combout\);

-- Location: FF_X60_Y3_N49
\RegFile[24][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[24][7]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][7]~q\);

-- Location: LABCELL_X62_Y4_N24
\Mux83~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux83~22_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[24][7]~q\))) # (\R.curInst\(15) & (\RegFile[25][7]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & (\RegFile[26][7]~q\)) # (\R.curInst\(15) & ((\RegFile[27][7]~q\)))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001110111011101110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[25][7]~q\,
	datac => \ALT_INV_RegFile[26][7]~q\,
	datad => \ALT_INV_RegFile[27][7]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][7]~q\,
	combout => \Mux83~22_combout\);

-- Location: LABCELL_X62_Y6_N36
\RegFile[28][7]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[28][7]~feeder_combout\ = ( \R.regWriteData\(7) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(7),
	combout => \RegFile[28][7]~feeder_combout\);

-- Location: FF_X62_Y6_N37
\RegFile[28][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[28][7]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][7]~q\);

-- Location: LABCELL_X62_Y4_N0
\Mux83~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux83~9_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux83~22_combout\)))) # (\R.curInst\(17) & ((!\Mux83~22_combout\ & ((\RegFile[28][7]~q\))) # (\Mux83~22_combout\ & (\RegFile[29][7]~q\))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) 
-- & (((\Mux83~22_combout\)))) # (\R.curInst\(17) & ((!\Mux83~22_combout\ & ((\RegFile[30][7]~DUPLICATE_q\))) # (\Mux83~22_combout\ & (\RegFile[31][7]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[29][7]~q\,
	datab => \ALT_INV_RegFile[31][7]~q\,
	datac => \ALT_INV_RegFile[30][7]~DUPLICATE_q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux83~22_combout\,
	datag => \ALT_INV_RegFile[28][7]~q\,
	combout => \Mux83~9_combout\);

-- Location: FF_X62_Y3_N44
\RegFile[3][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(7),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][7]~q\);

-- Location: FF_X68_Y7_N55
\RegFile[2][7]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[2][7]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][7]~DUPLICATE_q\);

-- Location: LABCELL_X60_Y3_N42
\RegFile[4][7]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[4][7]~feeder_combout\ = ( \R.regWriteData\(7) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(7),
	combout => \RegFile[4][7]~feeder_combout\);

-- Location: FF_X60_Y3_N43
\RegFile[4][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[4][7]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][7]~q\);

-- Location: LABCELL_X61_Y4_N3
\RegFile[6][7]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[6][7]~feeder_combout\ = ( \R.regWriteData\(7) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(7),
	combout => \RegFile[6][7]~feeder_combout\);

-- Location: FF_X61_Y4_N5
\RegFile[6][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[6][7]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][7]~q\);

-- Location: FF_X62_Y3_N14
\RegFile[5][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(7),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][7]~q\);

-- Location: FF_X62_Y3_N31
\RegFile[7][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(7),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][7]~q\);

-- Location: LABCELL_X62_Y3_N30
\Mux83~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux83~0_combout\ = ( \RegFile[7][7]~q\ & ( \R.curInst\(15) & ( (\RegFile[5][7]~q\) # (\R.curInst\(16)) ) ) ) # ( !\RegFile[7][7]~q\ & ( \R.curInst\(15) & ( (!\R.curInst\(16) & \RegFile[5][7]~q\) ) ) ) # ( \RegFile[7][7]~q\ & ( !\R.curInst\(15) & ( 
-- (!\R.curInst\(16) & (\RegFile[4][7]~q\)) # (\R.curInst\(16) & ((\RegFile[6][7]~q\))) ) ) ) # ( !\RegFile[7][7]~q\ & ( !\R.curInst\(15) & ( (!\R.curInst\(16) & (\RegFile[4][7]~q\)) # (\R.curInst\(16) & ((\RegFile[6][7]~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101001101010011010100110101001100000000111100000000111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[4][7]~q\,
	datab => \ALT_INV_RegFile[6][7]~q\,
	datac => \ALT_INV_R.curInst\(16),
	datad => \ALT_INV_RegFile[5][7]~q\,
	datae => \ALT_INV_RegFile[7][7]~q\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux83~0_combout\);

-- Location: MLABCELL_X59_Y7_N21
\RegFile[1][7]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[1][7]~feeder_combout\ = ( \R.regWriteData\(7) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(7),
	combout => \RegFile[1][7]~feeder_combout\);

-- Location: FF_X59_Y7_N22
\RegFile[1][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[1][7]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][7]~q\);

-- Location: LABCELL_X62_Y3_N42
\Mux83~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux83~26_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((\RegFile[1][7]~q\ & (\R.curInst\(15)))))) # (\R.curInst\(17) & ((((\Mux83~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & ((!\R.curInst\(15) & 
-- (((\RegFile[2][7]~DUPLICATE_q\)))) # (\R.curInst\(15) & (\RegFile[3][7]~q\)))) # (\R.curInst\(17) & ((((\Mux83~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001010000010100010001001010101010111110101111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[3][7]~q\,
	datac => \ALT_INV_RegFile[2][7]~DUPLICATE_q\,
	datad => \ALT_INV_R.curInst\(15),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux83~0_combout\,
	datag => \ALT_INV_RegFile[1][7]~q\,
	combout => \Mux83~26_combout\);

-- Location: FF_X68_Y7_N50
\RegFile[21][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(7),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][7]~q\);

-- Location: LABCELL_X64_Y4_N57
\RegFile[22][7]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[22][7]~feeder_combout\ = \R.regWriteData\(7)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.regWriteData\(7),
	combout => \RegFile[22][7]~feeder_combout\);

-- Location: FF_X64_Y4_N58
\RegFile[22][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[22][7]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][7]~q\);

-- Location: FF_X64_Y4_N44
\RegFile[23][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(7),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][7]~q\);

-- Location: FF_X63_Y5_N26
\RegFile[17][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(7),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][7]~q\);

-- Location: FF_X63_Y5_N2
\RegFile[18][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(7),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][7]~q\);

-- Location: FF_X64_Y4_N32
\RegFile[19][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(7),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][7]~q\);

-- Location: LABCELL_X63_Y5_N42
\RegFile[16][7]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[16][7]~feeder_combout\ = ( \R.regWriteData\(7) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(7),
	combout => \RegFile[16][7]~feeder_combout\);

-- Location: FF_X63_Y5_N44
\RegFile[16][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[16][7]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][7]~q\);

-- Location: LABCELL_X64_Y4_N30
\Mux83~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux83~18_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[16][7]~q\))) # (\R.curInst\(15) & (\RegFile[17][7]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & (\RegFile[18][7]~q\)) # (\R.curInst\(15) & ((\RegFile[19][7]~q\))))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[17][7]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[18][7]~q\,
	datad => \ALT_INV_RegFile[19][7]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][7]~q\,
	combout => \Mux83~18_combout\);

-- Location: FF_X59_Y4_N40
\RegFile[20][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(7),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][7]~q\);

-- Location: LABCELL_X64_Y4_N42
\Mux83~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux83~5_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux83~18_combout\))))) # (\R.curInst\(17) & (((!\Mux83~18_combout\ & ((\RegFile[20][7]~q\))) # (\Mux83~18_combout\ & (\RegFile[21][7]~q\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) 
-- & ((((\Mux83~18_combout\))))) # (\R.curInst\(17) & (((!\Mux83~18_combout\ & (\RegFile[22][7]~q\)) # (\Mux83~18_combout\ & ((\RegFile[23][7]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110111011101110111010101011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[21][7]~q\,
	datac => \ALT_INV_RegFile[22][7]~q\,
	datad => \ALT_INV_RegFile[23][7]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux83~18_combout\,
	datag => \ALT_INV_RegFile[20][7]~q\,
	combout => \Mux83~5_combout\);

-- Location: FF_X63_Y4_N20
\RegFile[15][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(7),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][7]~q\);

-- Location: FF_X61_Y7_N2
\RegFile[14][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(7),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][7]~q\);

-- Location: FF_X61_Y7_N26
\RegFile[13][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(7),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][7]~q\);

-- Location: FF_X64_Y3_N26
\RegFile[11][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(7),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][7]~q\);

-- Location: LABCELL_X64_Y3_N54
\RegFile[9][7]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[9][7]~feeder_combout\ = ( \R.regWriteData\(7) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(7),
	combout => \RegFile[9][7]~feeder_combout\);

-- Location: FF_X64_Y3_N55
\RegFile[9][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[9][7]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][7]~q\);

-- Location: FF_X64_Y3_N53
\RegFile[10][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(7),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][7]~q\);

-- Location: LABCELL_X66_Y5_N18
\RegFile[8][7]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[8][7]~feeder_combout\ = ( \R.regWriteData\(7) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(7),
	combout => \RegFile[8][7]~feeder_combout\);

-- Location: FF_X66_Y5_N19
\RegFile[8][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[8][7]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][7]~q\);

-- Location: LABCELL_X64_Y3_N24
\Mux83~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux83~14_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[8][7]~q\))) # (\R.curInst\(15) & (\RegFile[9][7]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[10][7]~q\))) # (\R.curInst\(15) & (\RegFile[11][7]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[11][7]~q\,
	datab => \ALT_INV_RegFile[9][7]~q\,
	datac => \ALT_INV_RegFile[10][7]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][7]~q\,
	combout => \Mux83~14_combout\);

-- Location: FF_X61_Y7_N43
\RegFile[12][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(7),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][7]~q\);

-- Location: LABCELL_X63_Y4_N18
\Mux83~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux83~1_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux83~14_combout\)))) # (\R.curInst\(17) & ((!\Mux83~14_combout\ & (\RegFile[12][7]~q\)) # (\Mux83~14_combout\ & ((\RegFile[13][7]~q\)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- ((((\Mux83~14_combout\))))) # (\R.curInst\(17) & (((!\Mux83~14_combout\ & ((\RegFile[14][7]~q\))) # (\Mux83~14_combout\ & (\RegFile[15][7]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111001100111111111101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][7]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[14][7]~q\,
	datad => \ALT_INV_RegFile[13][7]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux83~14_combout\,
	datag => \ALT_INV_RegFile[12][7]~q\,
	combout => \Mux83~1_combout\);

-- Location: LABCELL_X63_Y4_N39
\Mux83~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux83~13_combout\ = ( \Mux83~5_combout\ & ( \Mux83~1_combout\ & ( (!\R.curInst\(19) & (((\Mux83~26_combout\)) # (\R.curInst\(18)))) # (\R.curInst\(19) & ((!\R.curInst\(18)) # ((\Mux83~9_combout\)))) ) ) ) # ( !\Mux83~5_combout\ & ( \Mux83~1_combout\ & ( 
-- (!\R.curInst\(19) & (((\Mux83~26_combout\)) # (\R.curInst\(18)))) # (\R.curInst\(19) & (\R.curInst\(18) & (\Mux83~9_combout\))) ) ) ) # ( \Mux83~5_combout\ & ( !\Mux83~1_combout\ & ( (!\R.curInst\(19) & (!\R.curInst\(18) & ((\Mux83~26_combout\)))) # 
-- (\R.curInst\(19) & ((!\R.curInst\(18)) # ((\Mux83~9_combout\)))) ) ) ) # ( !\Mux83~5_combout\ & ( !\Mux83~1_combout\ & ( (!\R.curInst\(19) & (!\R.curInst\(18) & ((\Mux83~26_combout\)))) # (\R.curInst\(19) & (\R.curInst\(18) & (\Mux83~9_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000110001001010001011100110100100011101010110110011111101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(19),
	datab => \ALT_INV_R.curInst\(18),
	datac => \ALT_INV_Mux83~9_combout\,
	datad => \ALT_INV_Mux83~26_combout\,
	datae => \ALT_INV_Mux83~5_combout\,
	dataf => \ALT_INV_Mux83~1_combout\,
	combout => \Mux83~13_combout\);

-- Location: LABCELL_X74_Y7_N3
\Mux247~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux247~0_combout\ = ( \vAluSrc1~2_combout\ & ( (\R.curPC\(7) & !\vAluSrc1~1_combout\) ) ) # ( !\vAluSrc1~2_combout\ & ( (!\vAluSrc1~1_combout\ & \Mux83~13_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011110000000000001111000001010000010100000101000001010000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curPC\(7),
	datac => \ALT_INV_vAluSrc1~1_combout\,
	datad => \ALT_INV_Mux83~13_combout\,
	dataf => \ALT_INV_vAluSrc1~2_combout\,
	combout => \Mux247~0_combout\);

-- Location: FF_X74_Y7_N59
\Add2~25_OTERM723_NEW_REG828\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux247~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Add2~25_OTERM723_OTERM829\);

-- Location: LABCELL_X77_Y5_N24
\Mux148~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux148~0_combout\ = ( \R.curInst\(2) & ( \R.curInst\(26) & ( (!\R.curInst\(4) & (\R.curInst\(5) & \R.curInst\(6))) ) ) ) # ( !\R.curInst\(2) & ( \R.curInst\(26) & ( (!\R.curInst\(3) & ((!\R.curInst\(5) & ((!\R.curInst\(6)))) # (\R.curInst\(5) & 
-- (!\R.curInst\(4))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000010101000000010000000000000001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(3),
	datab => \ALT_INV_R.curInst\(4),
	datac => \ALT_INV_R.curInst\(5),
	datad => \ALT_INV_R.curInst\(6),
	datae => \ALT_INV_R.curInst\(2),
	dataf => \ALT_INV_R.curInst\(26),
	combout => \Mux148~0_combout\);

-- Location: LABCELL_X81_Y6_N12
\Add0~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~17_sumout\ = SUM(( \R.curPC\(6) ) + ( GND ) + ( \Add0~14\ ))
-- \Add0~18\ = CARRY(( \R.curPC\(6) ) + ( GND ) + ( \Add0~14\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.curPC\(6),
	cin => \Add0~14\,
	sumout => \Add0~17_sumout\,
	cout => \Add0~18\);

-- Location: LABCELL_X83_Y6_N27
\R.regWriteData[6]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.regWriteData[6]~feeder_combout\ = ( \Add0~17_sumout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_Add0~17_sumout\,
	combout => \R.regWriteData[6]~feeder_combout\);

-- Location: LABCELL_X74_Y7_N33
\Selector26~2_RTM0417\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector26~2_RTM0417_combout\ = ( \Mux248~0_combout\ & ( ((!\NxR.aluData2[6]~15_combout\ & (\R.aluOp.ALUOpXor_OTERM355\)) # (\NxR.aluData2[6]~15_combout\ & ((\R.aluOp.ALUOpAnd_OTERM357\)))) # (\R.aluOp.ALUOpOr_OTERM353\) ) ) # ( !\Mux248~0_combout\ & ( 
-- (\NxR.aluData2[6]~15_combout\ & ((\R.aluOp.ALUOpXor_OTERM355\) # (\R.aluOp.ALUOpOr_OTERM353\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000011100000111000001110000011101110101011111110111010101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpOr_OTERM353\,
	datab => \ALT_INV_R.aluOp.ALUOpXor_OTERM355\,
	datac => \ALT_INV_NxR.aluData2[6]~15_combout\,
	datad => \ALT_INV_R.aluOp.ALUOpAnd_OTERM357\,
	dataf => \ALT_INV_Mux248~0_combout\,
	combout => \Selector26~2_RTM0417_combout\);

-- Location: FF_X74_Y7_N34
\Selector26~2_NEW_REG414\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector26~2_RTM0417_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector26~2_OTERM415\);

-- Location: MLABCELL_X72_Y7_N33
\ShiftLeft0~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~2_combout\ = ( \NxR.aluData2[0]~16_combout\ & ( (\Mux253~0_combout\ & !\NxR.aluData2[1]~17_combout\) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (\Mux252~0_combout\)) # (\NxR.aluData2[1]~17_combout\ & 
-- ((\Mux254~0_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000110000111111000011000011111101000100010001000100010001000100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux253~0_combout\,
	datab => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datac => \ALT_INV_Mux252~0_combout\,
	datad => \ALT_INV_Mux254~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[0]~16_combout\,
	combout => \ShiftLeft0~2_combout\);

-- Location: FF_X72_Y7_N34
\ShiftLeft0~2_NEW_REG220\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~2_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~2_OTERM221\);

-- Location: LABCELL_X71_Y9_N45
\Selector27~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector27~0_combout\ = ( \R.aluOp.ALUOpSLL_OTERM359\ & ( !\NxR.aluData2[4]~20_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datae => \ALT_INV_R.aluOp.ALUOpSLL_OTERM359\,
	dataf => \ALT_INV_NxR.aluData2[4]~20_combout\,
	combout => \Selector27~0_combout\);

-- Location: FF_X71_Y9_N46
\Selector27~0_NEW_REG384\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector27~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector27~0_OTERM385\);

-- Location: FF_X64_Y5_N50
\RegFile[21][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(4),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][4]~q\);

-- Location: FF_X64_Y4_N56
\RegFile[22][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(4),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][4]~q\);

-- Location: FF_X63_Y5_N20
\RegFile[17][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(4),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][4]~q\);

-- Location: LABCELL_X63_Y5_N12
\RegFile[18][4]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[18][4]~feeder_combout\ = ( \R.regWriteData\(4) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(4),
	combout => \RegFile[18][4]~feeder_combout\);

-- Location: FF_X63_Y5_N13
\RegFile[18][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][4]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][4]~q\);

-- Location: FF_X63_Y7_N50
\RegFile[19][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(4),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][4]~q\);

-- Location: FF_X63_Y5_N38
\RegFile[16][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(4),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][4]~q\);

-- Location: LABCELL_X63_Y7_N48
\Mux86~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux86~18_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[16][4]~q\))) # (\R.curInst\(15) & (\RegFile[17][4]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & (\RegFile[18][4]~q\)) # (\R.curInst\(15) & ((\RegFile[19][4]~q\)))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001110111011101110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[17][4]~q\,
	datac => \ALT_INV_RegFile[18][4]~q\,
	datad => \ALT_INV_RegFile[19][4]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][4]~q\,
	combout => \Mux86~18_combout\);

-- Location: LABCELL_X56_Y7_N39
\RegFile[20][4]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[20][4]~feeder_combout\ = ( \R.regWriteData\(4) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(4),
	combout => \RegFile[20][4]~feeder_combout\);

-- Location: FF_X56_Y7_N40
\RegFile[20][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[20][4]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][4]~q\);

-- Location: LABCELL_X63_Y7_N21
\Mux86~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux86~5_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux86~18_combout\))))) # (\R.curInst\(17) & (((!\Mux86~18_combout\ & ((\RegFile[20][4]~q\))) # (\Mux86~18_combout\ & (\RegFile[21][4]~q\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) 
-- & ((((\Mux86~18_combout\))))) # (\R.curInst\(17) & (((!\Mux86~18_combout\ & (\RegFile[22][4]~q\)) # (\Mux86~18_combout\ & ((\RegFile[23][4]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110111011101110111010101011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[21][4]~q\,
	datac => \ALT_INV_RegFile[22][4]~q\,
	datad => \ALT_INV_RegFile[23][4]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux86~18_combout\,
	datag => \ALT_INV_RegFile[20][4]~q\,
	combout => \Mux86~5_combout\);

-- Location: FF_X62_Y7_N38
\RegFile[31][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(4),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][4]~q\);

-- Location: FF_X61_Y3_N44
\RegFile[29][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(4),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][4]~q\);

-- Location: LABCELL_X62_Y6_N54
\RegFile[30][4]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[30][4]~feeder_combout\ = ( \R.regWriteData\(4) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(4),
	combout => \RegFile[30][4]~feeder_combout\);

-- Location: FF_X62_Y6_N55
\RegFile[30][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[30][4]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][4]~q\);

-- Location: FF_X61_Y3_N50
\RegFile[25][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(4),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][4]~q\);

-- Location: FF_X61_Y3_N14
\RegFile[27][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(4),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][4]~q\);

-- Location: LABCELL_X53_Y3_N54
\RegFile[26][4]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[26][4]~feeder_combout\ = ( \R.regWriteData\(4) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(4),
	combout => \RegFile[26][4]~feeder_combout\);

-- Location: FF_X53_Y3_N55
\RegFile[26][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[26][4]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][4]~q\);

-- Location: LABCELL_X56_Y3_N3
\RegFile[24][4]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[24][4]~feeder_combout\ = ( \R.regWriteData\(4) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(4),
	combout => \RegFile[24][4]~feeder_combout\);

-- Location: FF_X56_Y3_N4
\RegFile[24][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[24][4]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][4]~q\);

-- Location: LABCELL_X61_Y3_N12
\Mux86~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux86~22_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[24][4]~q\))) # (\R.curInst\(15) & (\RegFile[25][4]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[26][4]~q\))) # (\R.curInst\(15) & (\RegFile[27][4]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[25][4]~q\,
	datab => \ALT_INV_RegFile[27][4]~q\,
	datac => \ALT_INV_RegFile[26][4]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][4]~q\,
	combout => \Mux86~22_combout\);

-- Location: LABCELL_X62_Y6_N48
\RegFile[28][4]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[28][4]~feeder_combout\ = ( \R.regWriteData\(4) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(4),
	combout => \RegFile[28][4]~feeder_combout\);

-- Location: FF_X62_Y6_N49
\RegFile[28][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[28][4]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][4]~q\);

-- Location: LABCELL_X62_Y7_N36
\Mux86~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux86~9_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux86~22_combout\)))) # (\R.curInst\(17) & ((!\Mux86~22_combout\ & ((\RegFile[28][4]~q\))) # (\Mux86~22_combout\ & (\RegFile[29][4]~q\))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) 
-- & (((\Mux86~22_combout\)))) # (\R.curInst\(17) & ((!\Mux86~22_combout\ & ((\RegFile[30][4]~q\))) # (\Mux86~22_combout\ & (\RegFile[31][4]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][4]~q\,
	datab => \ALT_INV_RegFile[29][4]~q\,
	datac => \ALT_INV_RegFile[30][4]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux86~22_combout\,
	datag => \ALT_INV_RegFile[28][4]~q\,
	combout => \Mux86~9_combout\);

-- Location: FF_X65_Y7_N2
\RegFile[2][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(4),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][4]~q\);

-- Location: LABCELL_X62_Y7_N54
\RegFile[3][4]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[3][4]~feeder_combout\ = ( \R.regWriteData\(4) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(4),
	combout => \RegFile[3][4]~feeder_combout\);

-- Location: FF_X62_Y7_N56
\RegFile[3][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[3][4]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][4]~q\);

-- Location: FF_X65_Y7_N31
\RegFile[5][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(4),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][4]~q\);

-- Location: LABCELL_X57_Y7_N6
\RegFile[6][4]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[6][4]~feeder_combout\ = ( \R.regWriteData\(4) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(4),
	combout => \RegFile[6][4]~feeder_combout\);

-- Location: FF_X57_Y7_N7
\RegFile[6][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[6][4]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][4]~q\);

-- Location: LABCELL_X60_Y3_N12
\RegFile[4][4]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[4][4]~feeder_combout\ = ( \R.regWriteData\(4) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(4),
	combout => \RegFile[4][4]~feeder_combout\);

-- Location: FF_X60_Y3_N13
\RegFile[4][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[4][4]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][4]~q\);

-- Location: FF_X65_Y7_N13
\RegFile[7][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(4),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][4]~q\);

-- Location: MLABCELL_X65_Y7_N12
\Mux86~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux86~0_combout\ = ( \RegFile[7][4]~q\ & ( \R.curInst\(15) & ( (\R.curInst\(16)) # (\RegFile[5][4]~q\) ) ) ) # ( !\RegFile[7][4]~q\ & ( \R.curInst\(15) & ( (\RegFile[5][4]~q\ & !\R.curInst\(16)) ) ) ) # ( \RegFile[7][4]~q\ & ( !\R.curInst\(15) & ( 
-- (!\R.curInst\(16) & ((\RegFile[4][4]~q\))) # (\R.curInst\(16) & (\RegFile[6][4]~q\)) ) ) ) # ( !\RegFile[7][4]~q\ & ( !\R.curInst\(15) & ( (!\R.curInst\(16) & ((\RegFile[4][4]~q\))) # (\R.curInst\(16) & (\RegFile[6][4]~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001111110011000000111111001101010000010100000101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[5][4]~q\,
	datab => \ALT_INV_RegFile[6][4]~q\,
	datac => \ALT_INV_R.curInst\(16),
	datad => \ALT_INV_RegFile[4][4]~q\,
	datae => \ALT_INV_RegFile[7][4]~q\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux86~0_combout\);

-- Location: MLABCELL_X59_Y7_N0
\RegFile[1][4]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[1][4]~feeder_combout\ = ( \R.regWriteData\(4) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(4),
	combout => \RegFile[1][4]~feeder_combout\);

-- Location: FF_X59_Y7_N2
\RegFile[1][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[1][4]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][4]~q\);

-- Location: LABCELL_X64_Y7_N42
\Mux86~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux86~26_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (\R.curInst\(15) & (\RegFile[1][4]~q\))) # (\R.curInst\(17) & ((((\Mux86~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & ((!\R.curInst\(15) & (\RegFile[2][4]~q\)) # 
-- (\R.curInst\(15) & (((\RegFile[3][4]~q\)))))) # (\R.curInst\(17) & ((((\Mux86~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010000000100000010000100110000110111001101110011101101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(15),
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[2][4]~q\,
	datad => \ALT_INV_RegFile[3][4]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux86~0_combout\,
	datag => \ALT_INV_RegFile[1][4]~q\,
	combout => \Mux86~26_combout\);

-- Location: FF_X64_Y5_N56
\RegFile[13][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(4),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][4]~q\);

-- Location: MLABCELL_X59_Y6_N24
\RegFile[14][4]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[14][4]~feeder_combout\ = ( \R.regWriteData\(4) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(4),
	combout => \RegFile[14][4]~feeder_combout\);

-- Location: FF_X59_Y6_N25
\RegFile[14][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[14][4]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][4]~q\);

-- Location: FF_X63_Y6_N14
\RegFile[15][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(4),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][4]~q\);

-- Location: FF_X63_Y6_N44
\RegFile[11][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(4),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][4]~q\);

-- Location: LABCELL_X64_Y3_N21
\RegFile[10][4]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[10][4]~feeder_combout\ = ( \R.regWriteData\(4) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(4),
	combout => \RegFile[10][4]~feeder_combout\);

-- Location: FF_X64_Y3_N22
\RegFile[10][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[10][4]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][4]~q\);

-- Location: FF_X64_Y5_N44
\RegFile[9][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(4),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][4]~q\);

-- Location: LABCELL_X63_Y6_N0
\RegFile[8][4]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[8][4]~feeder_combout\ = ( \R.regWriteData\(4) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(4),
	combout => \RegFile[8][4]~feeder_combout\);

-- Location: FF_X63_Y6_N1
\RegFile[8][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[8][4]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][4]~q\);

-- Location: LABCELL_X63_Y6_N42
\Mux86~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux86~14_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & (\RegFile[8][4]~q\)) # (\R.curInst\(15) & ((\RegFile[9][4]~q\)))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & ((\RegFile[10][4]~q\))) # (\R.curInst\(15) & (\RegFile[11][4]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001010101111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[11][4]~q\,
	datac => \ALT_INV_RegFile[10][4]~q\,
	datad => \ALT_INV_RegFile[9][4]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][4]~q\,
	combout => \Mux86~14_combout\);

-- Location: FF_X60_Y5_N4
\RegFile[12][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(4),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][4]~q\);

-- Location: LABCELL_X63_Y6_N12
\Mux86~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux86~1_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux86~14_combout\))))) # (\R.curInst\(17) & (((!\Mux86~14_combout\ & ((\RegFile[12][4]~q\))) # (\Mux86~14_combout\ & (\RegFile[13][4]~q\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) 
-- & ((((\Mux86~14_combout\))))) # (\R.curInst\(17) & (((!\Mux86~14_combout\ & (\RegFile[14][4]~q\)) # (\Mux86~14_combout\ & ((\RegFile[15][4]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110111011101110111010101011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[13][4]~q\,
	datac => \ALT_INV_RegFile[14][4]~q\,
	datad => \ALT_INV_RegFile[15][4]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux86~14_combout\,
	datag => \ALT_INV_RegFile[12][4]~q\,
	combout => \Mux86~1_combout\);

-- Location: LABCELL_X63_Y7_N42
\Mux86~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux86~13_combout\ = ( \Mux86~26_combout\ & ( \Mux86~1_combout\ & ( (!\R.curInst\(19)) # ((!\R.curInst\(18) & (\Mux86~5_combout\)) # (\R.curInst\(18) & ((\Mux86~9_combout\)))) ) ) ) # ( !\Mux86~26_combout\ & ( \Mux86~1_combout\ & ( (!\R.curInst\(18) & 
-- (\Mux86~5_combout\ & ((\R.curInst\(19))))) # (\R.curInst\(18) & (((!\R.curInst\(19)) # (\Mux86~9_combout\)))) ) ) ) # ( \Mux86~26_combout\ & ( !\Mux86~1_combout\ & ( (!\R.curInst\(18) & (((!\R.curInst\(19))) # (\Mux86~5_combout\))) # (\R.curInst\(18) & 
-- (((\Mux86~9_combout\ & \R.curInst\(19))))) ) ) ) # ( !\Mux86~26_combout\ & ( !\Mux86~1_combout\ & ( (\R.curInst\(19) & ((!\R.curInst\(18) & (\Mux86~5_combout\)) # (\R.curInst\(18) & ((\Mux86~9_combout\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001000111110011000100011100110011010001111111111101000111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux86~5_combout\,
	datab => \ALT_INV_R.curInst\(18),
	datac => \ALT_INV_Mux86~9_combout\,
	datad => \ALT_INV_R.curInst\(19),
	datae => \ALT_INV_Mux86~26_combout\,
	dataf => \ALT_INV_Mux86~1_combout\,
	combout => \Mux86~13_combout\);

-- Location: LABCELL_X73_Y7_N30
\Mux250~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux250~0_combout\ = ( !\vAluSrc1~1_combout\ & ( \Mux86~13_combout\ & ( (!\vAluSrc1~2_combout\) # (\R.curPC\(4)) ) ) ) # ( !\vAluSrc1~1_combout\ & ( !\Mux86~13_combout\ & ( (\R.curPC\(4) & \vAluSrc1~2_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000001111000000000000000011111111000011110000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.curPC\(4),
	datad => \ALT_INV_vAluSrc1~2_combout\,
	datae => \ALT_INV_vAluSrc1~1_combout\,
	dataf => \ALT_INV_Mux86~13_combout\,
	combout => \Mux250~0_combout\);

-- Location: LABCELL_X81_Y6_N0
\Add0~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~1_sumout\ = SUM(( \R.curPC\(2) ) + ( VCC ) + ( !VCC ))
-- \Add0~2\ = CARRY(( \R.curPC\(2) ) + ( VCC ) + ( !VCC ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.curPC\(2),
	cin => GND,
	sumout => \Add0~1_sumout\,
	cout => \Add0~2\);

-- Location: LABCELL_X81_Y6_N3
\Add0~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~5_sumout\ = SUM(( \R.curPC\(3) ) + ( GND ) + ( \Add0~2\ ))
-- \Add0~6\ = CARRY(( \R.curPC\(3) ) + ( GND ) + ( \Add0~2\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.curPC\(3),
	cin => \Add0~2\,
	sumout => \Add0~5_sumout\,
	cout => \Add0~6\);

-- Location: LABCELL_X81_Y6_N6
\Add0~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~9_sumout\ = SUM(( \R.curPC\(4) ) + ( GND ) + ( \Add0~6\ ))
-- \Add0~10\ = CARRY(( \R.curPC\(4) ) + ( GND ) + ( \Add0~6\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.curPC\(4),
	cin => \Add0~6\,
	sumout => \Add0~9_sumout\,
	cout => \Add0~10\);

-- Location: LABCELL_X81_Y6_N9
\Add0~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~13_sumout\ = SUM(( \R.curPC\(5) ) + ( GND ) + ( \Add0~10\ ))
-- \Add0~14\ = CARRY(( \R.curPC\(5) ) + ( GND ) + ( \Add0~10\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.curPC\(5),
	cin => \Add0~10\,
	sumout => \Add0~13_sumout\,
	cout => \Add0~14\);

-- Location: MLABCELL_X82_Y7_N6
\R.regWriteData[5]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.regWriteData[5]~feeder_combout\ = ( \Add0~13_sumout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_Add0~13_sumout\,
	combout => \R.regWriteData[5]~feeder_combout\);

-- Location: IOIBUF_X89_Y11_N61
\avm_d_readdata[29]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(29),
	o => \avm_d_readdata[29]~input_o\);

-- Location: LABCELL_X73_Y7_N24
\ShiftLeft0~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~7_combout\ = ( \NxR.aluData2[0]~16_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( \Mux252~0_combout\ ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( \Mux251~0_combout\ ) ) ) # ( \NxR.aluData2[0]~16_combout\ & ( 
-- !\NxR.aluData2[1]~17_combout\ & ( \Mux250~0_combout\ ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( !\NxR.aluData2[1]~17_combout\ & ( \Mux249~0_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101000000001111111100001111000011110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux249~0_combout\,
	datab => \ALT_INV_Mux252~0_combout\,
	datac => \ALT_INV_Mux251~0_combout\,
	datad => \ALT_INV_Mux250~0_combout\,
	datae => \ALT_INV_NxR.aluData2[0]~16_combout\,
	dataf => \ALT_INV_NxR.aluData2[1]~17_combout\,
	combout => \ShiftLeft0~7_combout\);

-- Location: FF_X73_Y7_N25
\ShiftLeft0~7_NEW_REG204\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~7_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~7_OTERM205\);

-- Location: LABCELL_X77_Y5_N27
\Mux149~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux149~1_combout\ = ( \R.curInst\(2) & ( \R.curInst\(25) & ( (!\R.curInst\(4) & (\R.curInst\(6) & \R.curInst\(5))) ) ) ) # ( !\R.curInst\(2) & ( \R.curInst\(25) & ( (!\R.curInst\(3) & ((!\R.curInst\(5) & ((!\R.curInst\(6)))) # (\R.curInst\(5) & 
-- (!\R.curInst\(4))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000010100000100010000000000000001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(3),
	datab => \ALT_INV_R.curInst\(4),
	datac => \ALT_INV_R.curInst\(6),
	datad => \ALT_INV_R.curInst\(5),
	datae => \ALT_INV_R.curInst\(2),
	dataf => \ALT_INV_R.curInst\(25),
	combout => \Mux149~1_combout\);

-- Location: FF_X66_Y7_N44
\RegFile[15][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(5),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][5]~q\);

-- Location: FF_X64_Y7_N50
\RegFile[13][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(5),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][5]~q\);

-- Location: LABCELL_X61_Y7_N57
\RegFile[14][5]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[14][5]~feeder_combout\ = ( \R.regWriteData\(5) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(5),
	combout => \RegFile[14][5]~feeder_combout\);

-- Location: FF_X61_Y7_N59
\RegFile[14][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[14][5]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][5]~q\);

-- Location: FF_X65_Y3_N38
\RegFile[11][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(5),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][5]~q\);

-- Location: MLABCELL_X65_Y3_N57
\RegFile[10][5]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[10][5]~feeder_combout\ = ( \R.regWriteData\(5) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(5),
	combout => \RegFile[10][5]~feeder_combout\);

-- Location: FF_X65_Y3_N58
\RegFile[10][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[10][5]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][5]~q\);

-- Location: FF_X65_Y3_N44
\RegFile[9][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(5),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][5]~q\);

-- Location: FF_X56_Y3_N19
\RegFile[8][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(5),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][5]~q\);

-- Location: MLABCELL_X65_Y3_N42
\Mux117~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux117~14_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & (\RegFile[8][5]~q\)) # (\R.curInst\(20) & ((\RegFile[9][5]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & ((\RegFile[10][5]~q\))) # (\R.curInst\(20) & (\RegFile[11][5]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110000110011111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[11][5]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[10][5]~q\,
	datad => \ALT_INV_RegFile[9][5]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][5]~q\,
	combout => \Mux117~14_combout\);

-- Location: FF_X66_Y7_N2
\RegFile[12][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(5),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][5]~q\);

-- Location: LABCELL_X64_Y7_N48
\Mux117~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux117~1_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux117~14_combout\)))) # (\R.curInst\(22) & ((!\Mux117~14_combout\ & ((\RegFile[12][5]~q\))) # (\Mux117~14_combout\ & (\RegFile[13][5]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux117~14_combout\)))) # (\R.curInst\(22) & ((!\Mux117~14_combout\ & ((\RegFile[14][5]~q\))) # (\Mux117~14_combout\ & (\RegFile[15][5]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][5]~q\,
	datab => \ALT_INV_RegFile[13][5]~q\,
	datac => \ALT_INV_RegFile[14][5]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux117~14_combout\,
	datag => \ALT_INV_RegFile[12][5]~q\,
	combout => \Mux117~1_combout\);

-- Location: FF_X62_Y7_N14
\RegFile[3][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(5),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][5]~q\);

-- Location: FF_X61_Y4_N41
\RegFile[2][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(5),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][5]~q\);

-- Location: LABCELL_X53_Y6_N51
\RegFile[4][5]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[4][5]~feeder_combout\ = ( \R.regWriteData\(5) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(5),
	combout => \RegFile[4][5]~feeder_combout\);

-- Location: FF_X53_Y6_N52
\RegFile[4][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[4][5]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][5]~q\);

-- Location: FF_X61_Y4_N17
\RegFile[7][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(5),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][5]~q\);

-- Location: FF_X60_Y3_N40
\RegFile[5][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(5),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][5]~q\);

-- Location: FF_X61_Y4_N31
\RegFile[6][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(5),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][5]~q\);

-- Location: LABCELL_X61_Y4_N51
\Mux117~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux117~0_combout\ = ( \R.curInst\(21) & ( \R.curInst\(20) & ( \RegFile[7][5]~q\ ) ) ) # ( !\R.curInst\(21) & ( \R.curInst\(20) & ( \RegFile[5][5]~q\ ) ) ) # ( \R.curInst\(21) & ( !\R.curInst\(20) & ( \RegFile[6][5]~q\ ) ) ) # ( !\R.curInst\(21) & ( 
-- !\R.curInst\(20) & ( \RegFile[4][5]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101000000001111111100001111000011110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[4][5]~q\,
	datab => \ALT_INV_RegFile[7][5]~q\,
	datac => \ALT_INV_RegFile[5][5]~q\,
	datad => \ALT_INV_RegFile[6][5]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	combout => \Mux117~0_combout\);

-- Location: MLABCELL_X59_Y7_N54
\RegFile[1][5]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[1][5]~feeder_combout\ = ( \R.regWriteData\(5) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(5),
	combout => \RegFile[1][5]~feeder_combout\);

-- Location: FF_X59_Y7_N55
\RegFile[1][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[1][5]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][5]~q\);

-- Location: LABCELL_X61_Y4_N39
\Mux117~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux117~26_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (\RegFile[1][5]~q\ & (\R.curInst\(20)))) # (\R.curInst\(22) & (((\Mux117~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (((\RegFile[2][5]~q\)))) # 
-- (\R.curInst\(20) & (\RegFile[3][5]~q\)))) # (\R.curInst\(22) & ((((\Mux117~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001100000011000100010000110011001111110011111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][5]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[2][5]~q\,
	datad => \ALT_INV_R.curInst\(20),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux117~0_combout\,
	datag => \ALT_INV_RegFile[1][5]~q\,
	combout => \Mux117~26_combout\);

-- Location: FF_X64_Y7_N23
\RegFile[21][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(5),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][5]~q\);

-- Location: LABCELL_X64_Y7_N54
\RegFile[23][5]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[23][5]~feeder_combout\ = ( \R.regWriteData\(5) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(5),
	combout => \RegFile[23][5]~feeder_combout\);

-- Location: FF_X64_Y7_N56
\RegFile[23][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[23][5]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][5]~q\);

-- Location: LABCELL_X56_Y7_N15
\RegFile[22][5]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[22][5]~feeder_combout\ = ( \R.regWriteData\(5) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(5),
	combout => \RegFile[22][5]~feeder_combout\);

-- Location: FF_X56_Y7_N16
\RegFile[22][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[22][5]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][5]~q\);

-- Location: FF_X63_Y7_N32
\RegFile[19][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(5),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][5]~q\);

-- Location: FF_X63_Y5_N16
\RegFile[18][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(5),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][5]~q\);

-- Location: FF_X63_Y7_N5
\RegFile[17][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(5),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][5]~q\);

-- Location: LABCELL_X60_Y7_N54
\RegFile[16][5]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[16][5]~feeder_combout\ = ( \R.regWriteData\(5) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(5),
	combout => \RegFile[16][5]~feeder_combout\);

-- Location: FF_X60_Y7_N55
\RegFile[16][5]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[16][5]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][5]~DUPLICATE_q\);

-- Location: LABCELL_X63_Y7_N3
\Mux117~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux117~18_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & (\RegFile[16][5]~DUPLICATE_q\)) # (\R.curInst\(20) & ((\RegFile[17][5]~q\)))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( 
-- (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[18][5]~q\))) # (\R.curInst\(20) & (\RegFile[19][5]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001010101111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[19][5]~q\,
	datac => \ALT_INV_RegFile[18][5]~q\,
	datad => \ALT_INV_RegFile[17][5]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][5]~DUPLICATE_q\,
	combout => \Mux117~18_combout\);

-- Location: LABCELL_X56_Y7_N9
\RegFile[20][5]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[20][5]~feeder_combout\ = ( \R.regWriteData\(5) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(5),
	combout => \RegFile[20][5]~feeder_combout\);

-- Location: FF_X56_Y7_N10
\RegFile[20][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[20][5]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][5]~q\);

-- Location: LABCELL_X64_Y7_N21
\Mux117~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux117~5_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux117~18_combout\)))) # (\R.curInst\(22) & ((!\Mux117~18_combout\ & ((\RegFile[20][5]~q\))) # (\Mux117~18_combout\ & (\RegFile[21][5]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux117~18_combout\)))) # (\R.curInst\(22) & ((!\Mux117~18_combout\ & ((\RegFile[22][5]~q\))) # (\Mux117~18_combout\ & (\RegFile[23][5]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][5]~q\,
	datab => \ALT_INV_RegFile[23][5]~q\,
	datac => \ALT_INV_RegFile[22][5]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux117~18_combout\,
	datag => \ALT_INV_RegFile[20][5]~q\,
	combout => \Mux117~5_combout\);

-- Location: FF_X62_Y7_N32
\RegFile[31][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(5),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][5]~q\);

-- Location: FF_X62_Y6_N47
\RegFile[30][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(5),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][5]~q\);

-- Location: LABCELL_X61_Y3_N36
\RegFile[27][5]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[27][5]~feeder_combout\ = ( \R.regWriteData\(5) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(5),
	combout => \RegFile[27][5]~feeder_combout\);

-- Location: FF_X61_Y3_N37
\RegFile[27][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[27][5]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][5]~q\);

-- Location: MLABCELL_X59_Y7_N36
\RegFile[25][5]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[25][5]~feeder_combout\ = ( \R.regWriteData\(5) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(5),
	combout => \RegFile[25][5]~feeder_combout\);

-- Location: FF_X59_Y7_N37
\RegFile[25][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[25][5]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][5]~q\);

-- Location: MLABCELL_X52_Y7_N21
\RegFile[26][5]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[26][5]~feeder_combout\ = ( \R.regWriteData\(5) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(5),
	combout => \RegFile[26][5]~feeder_combout\);

-- Location: FF_X52_Y7_N22
\RegFile[26][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[26][5]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][5]~q\);

-- Location: LABCELL_X64_Y6_N15
\RegFile[24][5]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[24][5]~feeder_combout\ = ( \R.regWriteData\(5) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(5),
	combout => \RegFile[24][5]~feeder_combout\);

-- Location: FF_X64_Y6_N16
\RegFile[24][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[24][5]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][5]~q\);

-- Location: LABCELL_X60_Y7_N33
\Mux117~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux117~22_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[24][5]~q\))) # (\R.curInst\(20) & (\RegFile[25][5]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[26][5]~q\))) # (\R.curInst\(20) & (\RegFile[27][5]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[27][5]~q\,
	datab => \ALT_INV_RegFile[25][5]~q\,
	datac => \ALT_INV_RegFile[26][5]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][5]~q\,
	combout => \Mux117~22_combout\);

-- Location: FF_X62_Y6_N26
\RegFile[28][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(5),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][5]~q\);

-- Location: LABCELL_X60_Y7_N18
\Mux117~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux117~9_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux117~22_combout\)))) # (\R.curInst\(22) & ((!\Mux117~22_combout\ & ((\RegFile[28][5]~q\))) # (\Mux117~22_combout\ & (\RegFile[29][5]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux117~22_combout\)))) # (\R.curInst\(22) & ((!\Mux117~22_combout\ & ((\RegFile[30][5]~q\))) # (\Mux117~22_combout\ & (\RegFile[31][5]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[29][5]~q\,
	datab => \ALT_INV_RegFile[31][5]~q\,
	datac => \ALT_INV_RegFile[30][5]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux117~22_combout\,
	datag => \ALT_INV_RegFile[28][5]~q\,
	combout => \Mux117~9_combout\);

-- Location: LABCELL_X64_Y7_N36
\Mux117~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux117~13_combout\ = ( \Mux117~5_combout\ & ( \Mux117~9_combout\ & ( ((!\R.curInst\(23) & ((\Mux117~26_combout\))) # (\R.curInst\(23) & (\Mux117~1_combout\))) # (\R.curInst\(24)) ) ) ) # ( !\Mux117~5_combout\ & ( \Mux117~9_combout\ & ( (!\R.curInst\(24) 
-- & ((!\R.curInst\(23) & ((\Mux117~26_combout\))) # (\R.curInst\(23) & (\Mux117~1_combout\)))) # (\R.curInst\(24) & (\R.curInst\(23))) ) ) ) # ( \Mux117~5_combout\ & ( !\Mux117~9_combout\ & ( (!\R.curInst\(24) & ((!\R.curInst\(23) & ((\Mux117~26_combout\))) 
-- # (\R.curInst\(23) & (\Mux117~1_combout\)))) # (\R.curInst\(24) & (!\R.curInst\(23))) ) ) ) # ( !\Mux117~5_combout\ & ( !\Mux117~9_combout\ & ( (!\R.curInst\(24) & ((!\R.curInst\(23) & ((\Mux117~26_combout\))) # (\R.curInst\(23) & (\Mux117~1_combout\)))) 
-- ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001010001010010001101100111000010011100110110101011111011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(24),
	datab => \ALT_INV_R.curInst\(23),
	datac => \ALT_INV_Mux117~1_combout\,
	datad => \ALT_INV_Mux117~26_combout\,
	datae => \ALT_INV_Mux117~5_combout\,
	dataf => \ALT_INV_Mux117~9_combout\,
	combout => \Mux117~13_combout\);

-- Location: MLABCELL_X72_Y5_N21
\NxR.aluData2[5]~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[5]~21_combout\ = ( \Mux117~13_combout\ & ( (!\vAluSrc2~1_combout\) # ((\Mux149~1_combout\ & \Equal4~1_combout\)) ) ) # ( !\Mux117~13_combout\ & ( (\Mux149~1_combout\ & (\vAluSrc2~1_combout\ & \Equal4~1_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000100000001000000010000000111001101110011011100110111001101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux149~1_combout\,
	datab => \ALT_INV_vAluSrc2~1_combout\,
	datac => \ALT_INV_Equal4~1_combout\,
	dataf => \ALT_INV_Mux117~13_combout\,
	combout => \NxR.aluData2[5]~21_combout\);

-- Location: MLABCELL_X72_Y5_N15
\Selector27~2_RTM0413\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector27~2_RTM0413_combout\ = ( \NxR.aluData2[5]~21_combout\ & ( ((!\Mux249~0_combout\ & (\R.aluOp.ALUOpXor_OTERM355\)) # (\Mux249~0_combout\ & ((\R.aluOp.ALUOpAnd_OTERM357\)))) # (\R.aluOp.ALUOpOr_OTERM353\) ) ) # ( !\NxR.aluData2[5]~21_combout\ & ( 
-- (\Mux249~0_combout\ & ((\R.aluOp.ALUOpXor_OTERM355\) # (\R.aluOp.ALUOpOr_OTERM353\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000011100000111000001110000011101110101011111110111010101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpOr_OTERM353\,
	datab => \ALT_INV_R.aluOp.ALUOpXor_OTERM355\,
	datac => \ALT_INV_Mux249~0_combout\,
	datad => \ALT_INV_R.aluOp.ALUOpAnd_OTERM357\,
	dataf => \ALT_INV_NxR.aluData2[5]~21_combout\,
	combout => \Selector27~2_RTM0413_combout\);

-- Location: FF_X72_Y5_N17
\Selector27~2_NEW_REG410\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector27~2_RTM0413_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector27~2_OTERM411\);

-- Location: MLABCELL_X72_Y7_N24
\ShiftLeft0~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~6_combout\ = ( \Mux254~0_combout\ & ( \Mux253~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (\NxR.aluData2[2]~19_combout\ & !\NxR.aluData2[3]~18_combout\)) ) ) ) # ( !\Mux254~0_combout\ & ( \Mux253~0_combout\ & ( 
-- (!\NxR.aluData2[0]~16_combout\ & (!\NxR.aluData2[1]~17_combout\ & (\NxR.aluData2[2]~19_combout\ & !\NxR.aluData2[3]~18_combout\))) ) ) ) # ( \Mux254~0_combout\ & ( !\Mux253~0_combout\ & ( (\NxR.aluData2[0]~16_combout\ & (!\NxR.aluData2[1]~17_combout\ & 
-- (\NxR.aluData2[2]~19_combout\ & !\NxR.aluData2[3]~18_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000001000000000000001000000000000000110000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datab => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datac => \ALT_INV_NxR.aluData2[2]~19_combout\,
	datad => \ALT_INV_NxR.aluData2[3]~18_combout\,
	datae => \ALT_INV_Mux254~0_combout\,
	dataf => \ALT_INV_Mux253~0_combout\,
	combout => \ShiftLeft0~6_combout\);

-- Location: FF_X72_Y7_N25
\ShiftLeft0~6_NEW_REG242\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~6_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~6_OTERM243\);

-- Location: LABCELL_X75_Y8_N45
\Selector27~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector27~3_combout\ = ( \ShiftLeft0~6_OTERM243\ & ( \ShiftRight0~7_OTERM233DUPLICATE_q\ & ( (!\Selector27~0_OTERM385\ & !\Selector27~2_OTERM411\) ) ) ) # ( !\ShiftLeft0~6_OTERM243\ & ( \ShiftRight0~7_OTERM233DUPLICATE_q\ & ( !\Selector27~2_OTERM411\ ) 
-- ) ) # ( \ShiftLeft0~6_OTERM243\ & ( !\ShiftRight0~7_OTERM233DUPLICATE_q\ & ( (!\Selector27~0_OTERM385\ & !\Selector27~2_OTERM411\) ) ) ) # ( !\ShiftLeft0~6_OTERM243\ & ( !\ShiftRight0~7_OTERM233DUPLICATE_q\ & ( (!\Selector27~2_OTERM411\ & 
-- ((!\ShiftLeft0~7_OTERM205\) # (!\Selector27~0_OTERM385\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1110000011100000110000001100000011110000111100001100000011000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~7_OTERM205\,
	datab => \ALT_INV_Selector27~0_OTERM385\,
	datac => \ALT_INV_Selector27~2_OTERM411\,
	datae => \ALT_INV_ShiftLeft0~6_OTERM243\,
	dataf => \ALT_INV_ShiftRight0~7_OTERM233DUPLICATE_q\,
	combout => \Selector27~3_combout\);

-- Location: LABCELL_X74_Y3_N12
\ShiftRight1~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~11_combout\ = ( \Mux230~0_combout\ & ( \NxR.aluData2[0]~16_combout\ & ( (\NxR.aluData2[1]~17_combout\) # (\Mux232~0_combout\) ) ) ) # ( !\Mux230~0_combout\ & ( \NxR.aluData2[0]~16_combout\ & ( (\Mux232~0_combout\ & 
-- !\NxR.aluData2[1]~17_combout\) ) ) ) # ( \Mux230~0_combout\ & ( !\NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((\Mux233~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux231~0_combout\)) ) ) ) # ( !\Mux230~0_combout\ & ( 
-- !\NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((\Mux233~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux231~0_combout\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100110011000011110011001101010101000000000101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux232~0_combout\,
	datab => \ALT_INV_Mux231~0_combout\,
	datac => \ALT_INV_Mux233~0_combout\,
	datad => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datae => \ALT_INV_Mux230~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[0]~16_combout\,
	combout => \ShiftRight1~11_combout\);

-- Location: FF_X74_Y3_N13
\ShiftRight1~11_NEW_REG34\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~11_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~11_OTERM35\);

-- Location: LABCELL_X74_Y8_N21
\ShiftRight0~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight0~8_combout\ = ( \ShiftRight0~0_OTERM17\ & ( (!\R.aluData2\(2) & (((\ShiftRight1~11_OTERM35\)) # (\R.aluData2\(3)))) # (\R.aluData2\(2) & (!\R.aluData2\(3) & (\ShiftRight1~12_OTERM57\))) ) ) # ( !\ShiftRight0~0_OTERM17\ & ( (!\R.aluData2\(3) & 
-- ((!\R.aluData2\(2) & ((\ShiftRight1~11_OTERM35\))) # (\R.aluData2\(2) & (\ShiftRight1~12_OTERM57\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010010001100000001001000110000100110101011100010011010101110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(2),
	datab => \ALT_INV_R.aluData2\(3),
	datac => \ALT_INV_ShiftRight1~12_OTERM57\,
	datad => \ALT_INV_ShiftRight1~11_OTERM35\,
	dataf => \ALT_INV_ShiftRight0~0_OTERM17\,
	combout => \ShiftRight0~8_combout\);

-- Location: LABCELL_X73_Y7_N18
\ShiftRight1~16\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~16_combout\ = ( \Mux247~0_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( (!\NxR.aluData2[0]~16_combout\) # (\Mux246~0_combout\) ) ) ) # ( !\Mux247~0_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( (\Mux246~0_combout\ & 
-- \NxR.aluData2[0]~16_combout\) ) ) ) # ( \Mux247~0_combout\ & ( !\NxR.aluData2[1]~17_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & ((\Mux249~0_combout\))) # (\NxR.aluData2[0]~16_combout\ & (\Mux248~0_combout\)) ) ) ) # ( !\Mux247~0_combout\ & ( 
-- !\NxR.aluData2[1]~17_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & ((\Mux249~0_combout\))) # (\NxR.aluData2[0]~16_combout\ & (\Mux248~0_combout\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001101010101001100110101010100000000000011111111111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux248~0_combout\,
	datab => \ALT_INV_Mux249~0_combout\,
	datac => \ALT_INV_Mux246~0_combout\,
	datad => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datae => \ALT_INV_Mux247~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[1]~17_combout\,
	combout => \ShiftRight1~16_combout\);

-- Location: FF_X73_Y7_N19
\ShiftRight1~16_NEW_REG208\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~16_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~16_OTERM209\);

-- Location: LABCELL_X75_Y7_N30
\ShiftRight1~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~17_combout\ = ( \Mux244~0_combout\ & ( \Mux243~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((\Mux245~0_combout\) # (\NxR.aluData2[0]~16_combout\)))) # (\NxR.aluData2[1]~17_combout\ & (((!\NxR.aluData2[0]~16_combout\)) # 
-- (\Mux242~0_combout\))) ) ) ) # ( !\Mux244~0_combout\ & ( \Mux243~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((!\NxR.aluData2[0]~16_combout\ & \Mux245~0_combout\)))) # (\NxR.aluData2[1]~17_combout\ & (((!\NxR.aluData2[0]~16_combout\)) # 
-- (\Mux242~0_combout\))) ) ) ) # ( \Mux244~0_combout\ & ( !\Mux243~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((\Mux245~0_combout\) # (\NxR.aluData2[0]~16_combout\)))) # (\NxR.aluData2[1]~17_combout\ & (\Mux242~0_combout\ & 
-- (\NxR.aluData2[0]~16_combout\))) ) ) ) # ( !\Mux244~0_combout\ & ( !\Mux243~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((!\NxR.aluData2[0]~16_combout\ & \Mux245~0_combout\)))) # (\NxR.aluData2[1]~17_combout\ & (\Mux242~0_combout\ & 
-- (\NxR.aluData2[0]~16_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000111000001000011011100110100110001111100010011110111111101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux242~0_combout\,
	datab => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datac => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datad => \ALT_INV_Mux245~0_combout\,
	datae => \ALT_INV_Mux244~0_combout\,
	dataf => \ALT_INV_Mux243~0_combout\,
	combout => \ShiftRight1~17_combout\);

-- Location: FF_X75_Y7_N31
\ShiftRight1~17_NEW_REG266\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~17_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~17_OTERM267\);

-- Location: FF_X61_Y2_N2
\RegFile[3][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(17),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][17]~q\);

-- Location: FF_X61_Y5_N8
\RegFile[2][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(17),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][17]~q\);

-- Location: LABCELL_X56_Y2_N45
\RegFile[4][17]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[4][17]~feeder_combout\ = ( \R.regWriteData\(17) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(17),
	combout => \RegFile[4][17]~feeder_combout\);

-- Location: FF_X56_Y2_N46
\RegFile[4][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[4][17]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][17]~q\);

-- Location: LABCELL_X61_Y4_N42
\RegFile[6][17]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[6][17]~feeder_combout\ = ( \R.regWriteData\(17) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(17),
	combout => \RegFile[6][17]~feeder_combout\);

-- Location: FF_X61_Y4_N43
\RegFile[6][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[6][17]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][17]~q\);

-- Location: FF_X61_Y2_N32
\RegFile[5][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(17),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][17]~q\);

-- Location: FF_X61_Y2_N25
\RegFile[7][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(17),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][17]~q\);

-- Location: LABCELL_X61_Y2_N24
\Mux73~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux73~0_combout\ = ( \RegFile[7][17]~q\ & ( \R.curInst\(15) & ( (\RegFile[5][17]~q\) # (\R.curInst\(16)) ) ) ) # ( !\RegFile[7][17]~q\ & ( \R.curInst\(15) & ( (!\R.curInst\(16) & \RegFile[5][17]~q\) ) ) ) # ( \RegFile[7][17]~q\ & ( !\R.curInst\(15) & ( 
-- (!\R.curInst\(16) & (\RegFile[4][17]~q\)) # (\R.curInst\(16) & ((\RegFile[6][17]~q\))) ) ) ) # ( !\RegFile[7][17]~q\ & ( !\R.curInst\(15) & ( (!\R.curInst\(16) & (\RegFile[4][17]~q\)) # (\R.curInst\(16) & ((\RegFile[6][17]~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010011100100111001001110010011100000000101010100101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(16),
	datab => \ALT_INV_RegFile[4][17]~q\,
	datac => \ALT_INV_RegFile[6][17]~q\,
	datad => \ALT_INV_RegFile[5][17]~q\,
	datae => \ALT_INV_RegFile[7][17]~q\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux73~0_combout\);

-- Location: FF_X61_Y5_N22
\RegFile[1][17]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(17),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][17]~DUPLICATE_q\);

-- Location: LABCELL_X61_Y2_N0
\Mux73~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux73~26_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (\RegFile[1][17]~DUPLICATE_q\ & (\R.curInst\(15)))) # (\R.curInst\(17) & (((\Mux73~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & ((!\R.curInst\(15) & 
-- (((\RegFile[2][17]~q\)))) # (\R.curInst\(15) & (\RegFile[3][17]~q\)))) # (\R.curInst\(17) & ((((\Mux73~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001100000011000100010000110011001111110011111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][17]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[2][17]~q\,
	datad => \ALT_INV_R.curInst\(15),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux73~0_combout\,
	datag => \ALT_INV_RegFile[1][17]~DUPLICATE_q\,
	combout => \Mux73~26_combout\);

-- Location: FF_X62_Y4_N56
\RegFile[31][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(17),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][17]~q\);

-- Location: FF_X66_Y3_N41
\RegFile[30][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(17),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][17]~q\);

-- Location: FF_X62_Y5_N44
\RegFile[29][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(17),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][17]~q\);

-- Location: FF_X62_Y4_N38
\RegFile[25][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(17),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][17]~q\);

-- Location: FF_X62_Y4_N20
\RegFile[27][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(17),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][17]~q\);

-- Location: LABCELL_X60_Y2_N15
\RegFile[26][17]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[26][17]~feeder_combout\ = ( \R.regWriteData\(17) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(17),
	combout => \RegFile[26][17]~feeder_combout\);

-- Location: FF_X60_Y2_N16
\RegFile[26][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[26][17]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][17]~q\);

-- Location: FF_X59_Y5_N34
\RegFile[24][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(17),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][17]~q\);

-- Location: LABCELL_X62_Y4_N18
\Mux73~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux73~22_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[24][17]~q\))) # (\R.curInst\(15) & (\RegFile[25][17]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[26][17]~q\))) # (\R.curInst\(15) & (\RegFile[27][17]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[25][17]~q\,
	datab => \ALT_INV_RegFile[27][17]~q\,
	datac => \ALT_INV_RegFile[26][17]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][17]~q\,
	combout => \Mux73~22_combout\);

-- Location: LABCELL_X60_Y6_N48
\RegFile[28][17]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[28][17]~feeder_combout\ = ( \R.regWriteData\(17) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(17),
	combout => \RegFile[28][17]~feeder_combout\);

-- Location: FF_X60_Y6_N49
\RegFile[28][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[28][17]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][17]~q\);

-- Location: LABCELL_X62_Y4_N54
\Mux73~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux73~9_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux73~22_combout\))))) # (\R.curInst\(17) & (((!\Mux73~22_combout\ & (\RegFile[28][17]~q\)) # (\Mux73~22_combout\ & ((\RegFile[29][17]~q\)))))) ) ) # ( \R.curInst\(16) & ( 
-- (!\R.curInst\(17) & ((((\Mux73~22_combout\))))) # (\R.curInst\(17) & (((!\Mux73~22_combout\ & ((\RegFile[30][17]~q\))) # (\Mux73~22_combout\ & (\RegFile[31][17]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110101010111111111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[31][17]~q\,
	datac => \ALT_INV_RegFile[30][17]~q\,
	datad => \ALT_INV_RegFile[29][17]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux73~22_combout\,
	datag => \ALT_INV_RegFile[28][17]~q\,
	combout => \Mux73~9_combout\);

-- Location: LABCELL_X62_Y5_N24
\RegFile[21][17]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[21][17]~feeder_combout\ = ( \R.regWriteData\(17) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(17),
	combout => \RegFile[21][17]~feeder_combout\);

-- Location: FF_X62_Y5_N25
\RegFile[21][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[21][17]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][17]~q\);

-- Location: FF_X63_Y4_N14
\RegFile[23][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(17),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][17]~q\);

-- Location: LABCELL_X61_Y6_N45
\RegFile[22][17]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[22][17]~feeder_combout\ = ( \R.regWriteData\(17) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(17),
	combout => \RegFile[22][17]~feeder_combout\);

-- Location: FF_X61_Y6_N46
\RegFile[22][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[22][17]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][17]~q\);

-- Location: FF_X63_Y5_N56
\RegFile[17][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(17),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][17]~q\);

-- Location: FF_X63_Y4_N44
\RegFile[19][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(17),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][17]~q\);

-- Location: LABCELL_X63_Y5_N6
\RegFile[18][17]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[18][17]~feeder_combout\ = \R.regWriteData\(17)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110011001100110011001100110011001100110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.regWriteData\(17),
	combout => \RegFile[18][17]~feeder_combout\);

-- Location: FF_X63_Y5_N7
\RegFile[18][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][17]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][17]~q\);

-- Location: LABCELL_X63_Y5_N36
\RegFile[16][17]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[16][17]~feeder_combout\ = ( \R.regWriteData\(17) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(17),
	combout => \RegFile[16][17]~feeder_combout\);

-- Location: FF_X63_Y5_N37
\RegFile[16][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[16][17]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][17]~q\);

-- Location: LABCELL_X63_Y4_N42
\Mux73~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux73~18_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[16][17]~q\))) # (\R.curInst\(15) & (\RegFile[17][17]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[18][17]~q\))) # (\R.curInst\(15) & (\RegFile[19][17]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[17][17]~q\,
	datab => \ALT_INV_RegFile[19][17]~q\,
	datac => \ALT_INV_RegFile[18][17]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][17]~q\,
	combout => \Mux73~18_combout\);

-- Location: FF_X59_Y5_N10
\RegFile[20][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(17),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][17]~q\);

-- Location: LABCELL_X63_Y4_N12
\Mux73~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux73~5_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux73~18_combout\)))) # (\R.curInst\(17) & ((!\Mux73~18_combout\ & ((\RegFile[20][17]~q\))) # (\Mux73~18_combout\ & (\RegFile[21][17]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux73~18_combout\)))) # (\R.curInst\(17) & ((!\Mux73~18_combout\ & ((\RegFile[22][17]~q\))) # (\Mux73~18_combout\ & (\RegFile[23][17]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][17]~q\,
	datab => \ALT_INV_RegFile[23][17]~q\,
	datac => \ALT_INV_RegFile[22][17]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux73~18_combout\,
	datag => \ALT_INV_RegFile[20][17]~q\,
	combout => \Mux73~5_combout\);

-- Location: FF_X63_Y4_N56
\RegFile[15][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(17),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][17]~q\);

-- Location: MLABCELL_X59_Y6_N57
\RegFile[14][17]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[14][17]~feeder_combout\ = ( \R.regWriteData\(17) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(17),
	combout => \RegFile[14][17]~feeder_combout\);

-- Location: FF_X59_Y6_N58
\RegFile[14][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[14][17]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][17]~q\);

-- Location: FF_X64_Y3_N2
\RegFile[11][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(17),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][17]~q\);

-- Location: FF_X64_Y3_N8
\RegFile[9][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(17),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][17]~q\);

-- Location: LABCELL_X64_Y3_N18
\RegFile[10][17]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[10][17]~feeder_combout\ = \R.regWriteData\(17)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.regWriteData\(17),
	combout => \RegFile[10][17]~feeder_combout\);

-- Location: FF_X64_Y3_N20
\RegFile[10][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[10][17]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][17]~q\);

-- Location: FF_X66_Y5_N8
\RegFile[8][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(17),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][17]~q\);

-- Location: LABCELL_X64_Y3_N0
\Mux73~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux73~14_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[8][17]~q\))) # (\R.curInst\(15) & (\RegFile[9][17]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[10][17]~q\))) # (\R.curInst\(15) & (\RegFile[11][17]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[11][17]~q\,
	datab => \ALT_INV_RegFile[9][17]~q\,
	datac => \ALT_INV_RegFile[10][17]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][17]~q\,
	combout => \Mux73~14_combout\);

-- Location: FF_X62_Y2_N7
\RegFile[12][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(17),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][17]~q\);

-- Location: LABCELL_X63_Y4_N54
\Mux73~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux73~1_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux73~14_combout\)))) # (\R.curInst\(17) & ((!\Mux73~14_combout\ & (\RegFile[12][17]~q\)) # (\Mux73~14_combout\ & ((\RegFile[13][17]~q\)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) 
-- & ((((\Mux73~14_combout\))))) # (\R.curInst\(17) & (((!\Mux73~14_combout\ & ((\RegFile[14][17]~q\))) # (\Mux73~14_combout\ & (\RegFile[15][17]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111001100111111111101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][17]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[14][17]~q\,
	datad => \ALT_INV_RegFile[13][17]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux73~14_combout\,
	datag => \ALT_INV_RegFile[12][17]~q\,
	combout => \Mux73~1_combout\);

-- Location: LABCELL_X62_Y4_N42
\Mux73~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux73~13_combout\ = ( \Mux73~5_combout\ & ( \Mux73~1_combout\ & ( (!\R.curInst\(18) & (((\R.curInst\(19))) # (\Mux73~26_combout\))) # (\R.curInst\(18) & (((!\R.curInst\(19)) # (\Mux73~9_combout\)))) ) ) ) # ( !\Mux73~5_combout\ & ( \Mux73~1_combout\ & ( 
-- (!\R.curInst\(18) & (\Mux73~26_combout\ & ((!\R.curInst\(19))))) # (\R.curInst\(18) & (((!\R.curInst\(19)) # (\Mux73~9_combout\)))) ) ) ) # ( \Mux73~5_combout\ & ( !\Mux73~1_combout\ & ( (!\R.curInst\(18) & (((\R.curInst\(19))) # (\Mux73~26_combout\))) # 
-- (\R.curInst\(18) & (((\Mux73~9_combout\ & \R.curInst\(19))))) ) ) ) # ( !\Mux73~5_combout\ & ( !\Mux73~1_combout\ & ( (!\R.curInst\(18) & (\Mux73~26_combout\ & ((!\R.curInst\(19))))) # (\R.curInst\(18) & (((\Mux73~9_combout\ & \R.curInst\(19))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010001000000101001000101010111101110111000001010111011110101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(18),
	datab => \ALT_INV_Mux73~26_combout\,
	datac => \ALT_INV_Mux73~9_combout\,
	datad => \ALT_INV_R.curInst\(19),
	datae => \ALT_INV_Mux73~5_combout\,
	dataf => \ALT_INV_Mux73~1_combout\,
	combout => \Mux73~13_combout\);

-- Location: LABCELL_X73_Y6_N0
\Mux237~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux237~0_combout\ = ( \Mux73~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC\(17)))) ) ) # ( !\Mux73~13_combout\ & ( (\vAluSrc1~2_combout\ & (\R.curPC\(17) & !\vAluSrc1~1_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000000000000110000000011001111000000001100111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_vAluSrc1~2_combout\,
	datac => \ALT_INV_R.curPC\(17),
	datad => \ALT_INV_vAluSrc1~1_combout\,
	dataf => \ALT_INV_Mux73~13_combout\,
	combout => \Mux237~0_combout\);

-- Location: LABCELL_X74_Y6_N42
\ShiftRight1~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~10_combout\ = ( \Mux234~0_combout\ & ( \Mux236~0_combout\ & ( ((!\NxR.aluData2[1]~17_combout\ & ((\Mux237~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux235~0_combout\))) # (\NxR.aluData2[0]~16_combout\) ) ) ) # ( !\Mux234~0_combout\ & 
-- ( \Mux236~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((\NxR.aluData2[0]~16_combout\) # (\Mux237~0_combout\)))) # (\NxR.aluData2[1]~17_combout\ & (\Mux235~0_combout\ & ((!\NxR.aluData2[0]~16_combout\)))) ) ) ) # ( \Mux234~0_combout\ & ( 
-- !\Mux236~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((\Mux237~0_combout\ & !\NxR.aluData2[0]~16_combout\)))) # (\NxR.aluData2[1]~17_combout\ & (((\NxR.aluData2[0]~16_combout\)) # (\Mux235~0_combout\))) ) ) ) # ( !\Mux234~0_combout\ & ( 
-- !\Mux236~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & ((!\NxR.aluData2[1]~17_combout\ & ((\Mux237~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux235~0_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001101100000000000110110101010100011011101010100001101111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datab => \ALT_INV_Mux235~0_combout\,
	datac => \ALT_INV_Mux237~0_combout\,
	datad => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datae => \ALT_INV_Mux234~0_combout\,
	dataf => \ALT_INV_Mux236~0_combout\,
	combout => \ShiftRight1~10_combout\);

-- Location: FF_X74_Y6_N43
\ShiftRight1~10_NEW_REG264\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~10_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~10_OTERM265\);

-- Location: MLABCELL_X78_Y9_N48
\ShiftRight1~42\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~42_combout\ = ( \ShiftRight1~17_OTERM267\ & ( \ShiftRight1~10_OTERM265\ & ( ((!\R.aluData2\(3) & (\ShiftRight1~16_OTERM209\)) # (\R.aluData2\(3) & ((\ShiftRight1~18_OTERM269\)))) # (\R.aluData2\(2)) ) ) ) # ( !\ShiftRight1~17_OTERM267\ & ( 
-- \ShiftRight1~10_OTERM265\ & ( (!\R.aluData2\(3) & (\ShiftRight1~16_OTERM209\ & ((!\R.aluData2\(2))))) # (\R.aluData2\(3) & (((\R.aluData2\(2)) # (\ShiftRight1~18_OTERM269\)))) ) ) ) # ( \ShiftRight1~17_OTERM267\ & ( !\ShiftRight1~10_OTERM265\ & ( 
-- (!\R.aluData2\(3) & (((\R.aluData2\(2))) # (\ShiftRight1~16_OTERM209\))) # (\R.aluData2\(3) & (((\ShiftRight1~18_OTERM269\ & !\R.aluData2\(2))))) ) ) ) # ( !\ShiftRight1~17_OTERM267\ & ( !\ShiftRight1~10_OTERM265\ & ( (!\R.aluData2\(2) & 
-- ((!\R.aluData2\(3) & (\ShiftRight1~16_OTERM209\)) # (\R.aluData2\(3) & ((\ShiftRight1~18_OTERM269\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100011100000000010001111100110001000111001100110100011111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~16_OTERM209\,
	datab => \ALT_INV_R.aluData2\(3),
	datac => \ALT_INV_ShiftRight1~18_OTERM269\,
	datad => \ALT_INV_R.aluData2\(2),
	datae => \ALT_INV_ShiftRight1~17_OTERM267\,
	dataf => \ALT_INV_ShiftRight1~10_OTERM265\,
	combout => \ShiftRight1~42_combout\);

-- Location: LABCELL_X75_Y8_N51
\Selector27~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector27~4_combout\ = ( \ShiftRight0~8_combout\ & ( \ShiftRight1~42_combout\ & ( (!\Selector31~5_OTERM599\ & (\Selector27~3_combout\ & !\Selector31~7_OTERM383\)) ) ) ) # ( !\ShiftRight0~8_combout\ & ( \ShiftRight1~42_combout\ & ( 
-- (!\Selector31~5_OTERM599\ & \Selector27~3_combout\) ) ) ) # ( \ShiftRight0~8_combout\ & ( !\ShiftRight1~42_combout\ & ( (\Selector27~3_combout\ & !\Selector31~7_OTERM383\) ) ) ) # ( !\ShiftRight0~8_combout\ & ( !\ShiftRight1~42_combout\ & ( 
-- \Selector27~3_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110011001100000011000000100010001000100010000000100000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector31~5_OTERM599\,
	datab => \ALT_INV_Selector27~3_combout\,
	datac => \ALT_INV_Selector31~7_OTERM383\,
	datae => \ALT_INV_ShiftRight0~8_combout\,
	dataf => \ALT_INV_ShiftRight1~42_combout\,
	combout => \Selector27~4_combout\);

-- Location: FF_X72_Y5_N47
\Add2~17_OTERM727_NEW_REG840\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \NxR.aluData2[5]~21_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Add2~17_OTERM727_OTERM841\);

-- Location: FF_X78_Y6_N17
\R.aluData1[5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux249~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData1\(5));

-- Location: FF_X73_Y7_N10
\R.aluData1[4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux250~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData1\(4));

-- Location: FF_X72_Y7_N46
\R.aluData1[3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux251~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData1\(3));

-- Location: FF_X72_Y7_N52
\R.aluData1[2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux252~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData1\(2));

-- Location: MLABCELL_X78_Y6_N6
\Add1~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~9_sumout\ = SUM(( \R.aluData2\(2) ) + ( \R.aluData1\(2) ) + ( \Add1~6\ ))
-- \Add1~10\ = CARRY(( \R.aluData2\(2) ) + ( \R.aluData1\(2) ) + ( \Add1~6\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluData1\(2),
	datad => \ALT_INV_R.aluData2\(2),
	cin => \Add1~6\,
	sumout => \Add1~9_sumout\,
	cout => \Add1~10\);

-- Location: MLABCELL_X78_Y6_N9
\Add1~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~13_sumout\ = SUM(( \R.aluData1\(3) ) + ( \R.aluData2\(3) ) + ( \Add1~10\ ))
-- \Add1~14\ = CARRY(( \R.aluData1\(3) ) + ( \R.aluData2\(3) ) + ( \Add1~10\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluData2\(3),
	datad => \ALT_INV_R.aluData1\(3),
	cin => \Add1~10\,
	sumout => \Add1~13_sumout\,
	cout => \Add1~14\);

-- Location: MLABCELL_X78_Y6_N12
\Add1~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~17_sumout\ = SUM(( \R.aluData1\(4) ) + ( \R.aluData2\(4) ) + ( \Add1~14\ ))
-- \Add1~18\ = CARRY(( \R.aluData1\(4) ) + ( \R.aluData2\(4) ) + ( \Add1~14\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluData2\(4),
	datad => \ALT_INV_R.aluData1\(4),
	cin => \Add1~14\,
	sumout => \Add1~17_sumout\,
	cout => \Add1~18\);

-- Location: MLABCELL_X78_Y6_N15
\Add1~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~21_sumout\ = SUM(( \Add2~17_OTERM727_OTERM841\ ) + ( \R.aluData1\(5) ) + ( \Add1~18\ ))
-- \Add1~22\ = CARRY(( \Add2~17_OTERM727_OTERM841\ ) + ( \R.aluData1\(5) ) + ( \Add1~18\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add2~17_OTERM727_OTERM841\,
	datac => \ALT_INV_R.aluData1\(5),
	cin => \Add1~18\,
	sumout => \Add1~21_sumout\,
	cout => \Add1~22\);

-- Location: LABCELL_X79_Y6_N6
\Add2~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~9_sumout\ = SUM(( !\R.aluData1\(2) $ (\R.aluData2\(2)) ) + ( \Add2~7\ ) + ( \Add2~6\ ))
-- \Add2~10\ = CARRY(( !\R.aluData1\(2) $ (\R.aluData2\(2)) ) + ( \Add2~7\ ) + ( \Add2~6\ ))
-- \Add2~11\ = SHARE((\R.aluData1\(2) & !\R.aluData2\(2)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000000000000000000000001111000000001111",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluData1\(2),
	datad => \ALT_INV_R.aluData2\(2),
	cin => \Add2~6\,
	sharein => \Add2~7\,
	sumout => \Add2~9_sumout\,
	cout => \Add2~10\,
	shareout => \Add2~11\);

-- Location: LABCELL_X79_Y6_N9
\Add2~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~13_sumout\ = SUM(( !\R.aluData2\(3) $ (\R.aluData1\(3)) ) + ( \Add2~11\ ) + ( \Add2~10\ ))
-- \Add2~14\ = CARRY(( !\R.aluData2\(3) $ (\R.aluData1\(3)) ) + ( \Add2~11\ ) + ( \Add2~10\ ))
-- \Add2~15\ = SHARE((!\R.aluData2\(3) & \R.aluData1\(3)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000001111000000000000000000001111000000001111",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluData2\(3),
	datad => \ALT_INV_R.aluData1\(3),
	cin => \Add2~10\,
	sharein => \Add2~11\,
	sumout => \Add2~13_sumout\,
	cout => \Add2~14\,
	shareout => \Add2~15\);

-- Location: LABCELL_X79_Y6_N12
\Add2~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~17_sumout\ = SUM(( !\R.aluData1\(4) $ (\R.aluData2\(4)) ) + ( \Add2~15\ ) + ( \Add2~14\ ))
-- \Add2~18\ = CARRY(( !\R.aluData1\(4) $ (\R.aluData2\(4)) ) + ( \Add2~15\ ) + ( \Add2~14\ ))
-- \Add2~19\ = SHARE((\R.aluData1\(4) & !\R.aluData2\(4)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000000000000000000000001111000000001111",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluData1\(4),
	datad => \ALT_INV_R.aluData2\(4),
	cin => \Add2~14\,
	sharein => \Add2~15\,
	sumout => \Add2~17_sumout\,
	cout => \Add2~18\,
	shareout => \Add2~19\);

-- Location: LABCELL_X79_Y6_N15
\Add2~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~21_sumout\ = SUM(( !\Add2~17_OTERM727_OTERM841\ $ (\R.aluData1\(5)) ) + ( \Add2~19\ ) + ( \Add2~18\ ))
-- \Add2~22\ = CARRY(( !\Add2~17_OTERM727_OTERM841\ $ (\R.aluData1\(5)) ) + ( \Add2~19\ ) + ( \Add2~18\ ))
-- \Add2~23\ = SHARE((!\Add2~17_OTERM727_OTERM841\ & \R.aluData1\(5)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000010100000101000000000000000001010010110100101",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add2~17_OTERM727_OTERM841\,
	datac => \ALT_INV_R.aluData1\(5),
	cin => \Add2~18\,
	sharein => \Add2~19\,
	sumout => \Add2~21_sumout\,
	cout => \Add2~22\,
	shareout => \Add2~23\);

-- Location: MLABCELL_X82_Y7_N45
\Selector27~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector27~1_combout\ = ( \Add2~21_sumout\ & ( ((\R.aluOp.ALUOpAdd~q\ & \Add1~21_sumout\)) # (\R.aluOp.ALUOpSub~q\) ) ) # ( !\Add2~21_sumout\ & ( (\R.aluOp.ALUOpAdd~q\ & \Add1~21_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000001111000000000000111101010101010111110101010101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_Add1~21_sumout\,
	dataf => \ALT_INV_Add2~21_sumout\,
	combout => \Selector27~1_combout\);

-- Location: MLABCELL_X82_Y7_N30
\Comb:vRegWriteData[5]~0_RESYN1092\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[5]~0_RESYN1092_BDD1093\ = ( \ShiftRight1~41_combout\ & ( \Mux222~0_combout\ & ( ((!\R.aluCalc~q\ & ((\R.aluRes\(5)))) # (\R.aluCalc~q\ & (\Selector31~6_OTERM381\))) # (\R.memToReg~q\) ) ) ) # ( !\ShiftRight1~41_combout\ & ( 
-- \Mux222~0_combout\ & ( ((!\R.aluCalc~q\ & \R.aluRes\(5))) # (\R.memToReg~q\) ) ) ) # ( \ShiftRight1~41_combout\ & ( !\Mux222~0_combout\ & ( (!\R.memToReg~q\ & ((!\R.aluCalc~q\ & ((\R.aluRes\(5)))) # (\R.aluCalc~q\ & (\Selector31~6_OTERM381\)))) ) ) ) # ( 
-- !\ShiftRight1~41_combout\ & ( !\Mux222~0_combout\ & ( (!\R.aluCalc~q\ & (!\R.memToReg~q\ & \R.aluRes\(5))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011000000000100001101000000001111110011110001111111011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector31~6_OTERM381\,
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_R.memToReg~q\,
	datad => \ALT_INV_R.aluRes\(5),
	datae => \ALT_INV_ShiftRight1~41_combout\,
	dataf => \ALT_INV_Mux222~0_combout\,
	combout => \Comb:vRegWriteData[5]~0_RESYN1092_BDD1093\);

-- Location: MLABCELL_X82_Y7_N48
\Comb:vRegWriteData[5]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[5]~0_combout\ = ( \Selector27~1_combout\ & ( \Comb:vRegWriteData[5]~0_RESYN1092_BDD1093\ & ( (!\R.memToReg~q\) # (\avm_d_readdata[29]~input_o\) ) ) ) # ( !\Selector27~1_combout\ & ( \Comb:vRegWriteData[5]~0_RESYN1092_BDD1093\ & ( 
-- (!\R.memToReg~q\) # (\avm_d_readdata[29]~input_o\) ) ) ) # ( \Selector27~1_combout\ & ( !\Comb:vRegWriteData[5]~0_RESYN1092_BDD1093\ & ( (\R.aluCalc~q\ & !\R.memToReg~q\) ) ) ) # ( !\Selector27~1_combout\ & ( !\Comb:vRegWriteData[5]~0_RESYN1092_BDD1093\ & 
-- ( (\R.aluCalc~q\ & (!\R.memToReg~q\ & !\Selector27~4_combout\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011000000000000001100000011000011110101111101011111010111110101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_avm_d_readdata[29]~input_o\,
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_R.memToReg~q\,
	datad => \ALT_INV_Selector27~4_combout\,
	datae => \ALT_INV_Selector27~1_combout\,
	dataf => \ALT_INV_Comb:vRegWriteData[5]~0_RESYN1092_BDD1093\,
	combout => \Comb:vRegWriteData[5]~0_combout\);

-- Location: LABCELL_X71_Y7_N0
\Selector16~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector16~0_combout\ = ( \R.aluOp.ALUOpSLL_OTERM359\ & ( (\NxR.aluData2[4]~20_combout\ & (!\NxR.aluData2[2]~19_combout\ & !\NxR.aluData2[3]~18_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000110000000000000011000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_NxR.aluData2[4]~20_combout\,
	datac => \ALT_INV_NxR.aluData2[2]~19_combout\,
	datad => \ALT_INV_NxR.aluData2[3]~18_combout\,
	dataf => \ALT_INV_R.aluOp.ALUOpSLL_OTERM359\,
	combout => \Selector16~0_combout\);

-- Location: FF_X71_Y7_N1
\Selector16~0_NEW_REG392\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector16~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector16~0_OTERM393\);

-- Location: LABCELL_X75_Y4_N45
\Mux135~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux135~0_combout\ = ( \Mux123~2_combout\ & ( \R.curInst\(19) ) ) # ( !\Mux123~2_combout\ & ( \R.curInst\(19) & ( ((\vAluSrc1~0_combout\ & ((\R.curInst\(2)) # (\Mux124~0_combout\)))) # (\Mux149~0_combout\) ) ) ) # ( \Mux123~2_combout\ & ( !\R.curInst\(19) 
-- ) ) # ( !\Mux123~2_combout\ & ( !\R.curInst\(19) & ( (\Mux124~0_combout\ & \vAluSrc1~0_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101111111111111111100000111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux124~0_combout\,
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_vAluSrc1~0_combout\,
	datad => \ALT_INV_Mux149~0_combout\,
	datae => \ALT_INV_Mux123~2_combout\,
	dataf => \ALT_INV_R.curInst\(19),
	combout => \Mux135~0_combout\);

-- Location: FF_X72_Y1_N38
\RegFile[23][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(19),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][19]~q\);

-- Location: FF_X71_Y1_N38
\RegFile[21][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(19),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][19]~q\);

-- Location: LABCELL_X71_Y1_N21
\RegFile[22][19]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[22][19]~feeder_combout\ = ( \R.regWriteData\(19) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(19),
	combout => \RegFile[22][19]~feeder_combout\);

-- Location: FF_X71_Y1_N23
\RegFile[22][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[22][19]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][19]~q\);

-- Location: FF_X72_Y1_N50
\RegFile[19][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(19),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][19]~q\);

-- Location: FF_X72_Y1_N32
\RegFile[17][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(19),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][19]~q\);

-- Location: MLABCELL_X59_Y1_N36
\RegFile[18][19]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[18][19]~feeder_combout\ = ( \R.regWriteData\(19) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(19),
	combout => \RegFile[18][19]~feeder_combout\);

-- Location: FF_X59_Y1_N37
\RegFile[18][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][19]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][19]~q\);

-- Location: FF_X64_Y1_N2
\RegFile[16][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(19),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][19]~q\);

-- Location: MLABCELL_X72_Y1_N30
\Mux103~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux103~18_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[16][19]~q\))) # (\R.curInst\(20) & (\RegFile[17][19]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[18][19]~q\))) # (\R.curInst\(20) & (\RegFile[19][19]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[19][19]~q\,
	datab => \ALT_INV_RegFile[17][19]~q\,
	datac => \ALT_INV_RegFile[18][19]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][19]~q\,
	combout => \Mux103~18_combout\);

-- Location: FF_X74_Y1_N58
\RegFile[20][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(19),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][19]~q\);

-- Location: LABCELL_X71_Y1_N36
\Mux103~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux103~5_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux103~18_combout\)))) # (\R.curInst\(22) & ((!\Mux103~18_combout\ & ((\RegFile[20][19]~q\))) # (\Mux103~18_combout\ & (\RegFile[21][19]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux103~18_combout\)))) # (\R.curInst\(22) & ((!\Mux103~18_combout\ & ((\RegFile[22][19]~q\))) # (\Mux103~18_combout\ & (\RegFile[23][19]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[23][19]~q\,
	datab => \ALT_INV_RegFile[21][19]~q\,
	datac => \ALT_INV_RegFile[22][19]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux103~18_combout\,
	datag => \ALT_INV_RegFile[20][19]~q\,
	combout => \Mux103~5_combout\);

-- Location: FF_X72_Y3_N8
\RegFile[2][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(19),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][19]~q\);

-- Location: FF_X73_Y3_N49
\RegFile[7][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(19),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][19]~q\);

-- Location: LABCELL_X71_Y3_N27
\RegFile[6][19]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[6][19]~feeder_combout\ = ( \R.regWriteData\(19) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(19),
	combout => \RegFile[6][19]~feeder_combout\);

-- Location: FF_X71_Y3_N28
\RegFile[6][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[6][19]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][19]~q\);

-- Location: FF_X67_Y5_N47
\RegFile[4][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(19),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][19]~q\);

-- Location: FF_X72_Y3_N26
\RegFile[5][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(19),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][19]~q\);

-- Location: MLABCELL_X72_Y3_N24
\Mux103~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux103~0_combout\ = ( \RegFile[5][19]~q\ & ( \R.curInst\(20) & ( (!\R.curInst\(21)) # (\RegFile[7][19]~q\) ) ) ) # ( !\RegFile[5][19]~q\ & ( \R.curInst\(20) & ( (\RegFile[7][19]~q\ & \R.curInst\(21)) ) ) ) # ( \RegFile[5][19]~q\ & ( !\R.curInst\(20) & ( 
-- (!\R.curInst\(21) & ((\RegFile[4][19]~q\))) # (\R.curInst\(21) & (\RegFile[6][19]~q\)) ) ) ) # ( !\RegFile[5][19]~q\ & ( !\R.curInst\(20) & ( (!\R.curInst\(21) & ((\RegFile[4][19]~q\))) # (\R.curInst\(21) & (\RegFile[6][19]~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001111110011000000111111001100000101000001011111010111110101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[7][19]~q\,
	datab => \ALT_INV_RegFile[6][19]~q\,
	datac => \ALT_INV_R.curInst\(21),
	datad => \ALT_INV_RegFile[4][19]~q\,
	datae => \ALT_INV_RegFile[5][19]~q\,
	dataf => \ALT_INV_R.curInst\(20),
	combout => \Mux103~0_combout\);

-- Location: MLABCELL_X72_Y3_N57
\RegFile[1][19]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[1][19]~feeder_combout\ = ( \R.regWriteData\(19) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(19),
	combout => \RegFile[1][19]~feeder_combout\);

-- Location: FF_X72_Y3_N59
\RegFile[1][19]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[1][19]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][19]~DUPLICATE_q\);

-- Location: MLABCELL_X72_Y3_N6
\Mux103~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux103~26_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((\RegFile[1][19]~DUPLICATE_q\ & (\R.curInst\(20)))))) # (\R.curInst\(22) & ((((\Mux103~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & 
-- (((\RegFile[2][19]~q\)))) # (\R.curInst\(20) & (\RegFile[3][19]~q\)))) # (\R.curInst\(22) & ((((\Mux103~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001010000010100010001001010101010111110101111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[3][19]~q\,
	datac => \ALT_INV_RegFile[2][19]~q\,
	datad => \ALT_INV_R.curInst\(20),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux103~0_combout\,
	datag => \ALT_INV_RegFile[1][19]~DUPLICATE_q\,
	combout => \Mux103~26_combout\);

-- Location: FF_X66_Y2_N44
\RegFile[29][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(19),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][19]~q\);

-- Location: FF_X66_Y3_N47
\RegFile[30][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(19),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][19]~q\);

-- Location: FF_X66_Y3_N14
\RegFile[31][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(19),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][19]~q\);

-- Location: FF_X66_Y2_N20
\RegFile[25][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(19),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][19]~q\);

-- Location: FF_X66_Y2_N8
\RegFile[27][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(19),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][19]~q\);

-- Location: LABCELL_X60_Y2_N21
\RegFile[26][19]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[26][19]~feeder_combout\ = ( \R.regWriteData\(19) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(19),
	combout => \RegFile[26][19]~feeder_combout\);

-- Location: FF_X60_Y2_N22
\RegFile[26][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[26][19]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][19]~q\);

-- Location: FF_X59_Y2_N25
\RegFile[24][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(19),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][19]~q\);

-- Location: LABCELL_X66_Y2_N18
\Mux103~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux103~22_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[24][19]~q\))) # (\R.curInst\(20) & (\RegFile[25][19]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[26][19]~q\))) # (\R.curInst\(20) & (\RegFile[27][19]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[25][19]~q\,
	datab => \ALT_INV_RegFile[27][19]~q\,
	datac => \ALT_INV_RegFile[26][19]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][19]~q\,
	combout => \Mux103~22_combout\);

-- Location: FF_X66_Y3_N20
\RegFile[28][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(19),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][19]~q\);

-- Location: LABCELL_X66_Y2_N42
\Mux103~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux103~9_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux103~22_combout\))))) # (\R.curInst\(22) & (((!\Mux103~22_combout\ & ((\RegFile[28][19]~q\))) # (\Mux103~22_combout\ & (\RegFile[29][19]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- (!\R.curInst\(22) & ((((\Mux103~22_combout\))))) # (\R.curInst\(22) & (((!\Mux103~22_combout\ & (\RegFile[30][19]~q\)) # (\Mux103~22_combout\ & ((\RegFile[31][19]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110111011101110111010101011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[29][19]~q\,
	datac => \ALT_INV_RegFile[30][19]~q\,
	datad => \ALT_INV_RegFile[31][19]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux103~22_combout\,
	datag => \ALT_INV_RegFile[28][19]~q\,
	combout => \Mux103~9_combout\);

-- Location: FF_X63_Y1_N56
\RegFile[13][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(19),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][19]~q\);

-- Location: FF_X63_Y3_N56
\RegFile[15][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(19),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][19]~q\);

-- Location: FF_X63_Y3_N53
\RegFile[14][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(19),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][19]~q\);

-- Location: FF_X63_Y1_N2
\RegFile[9][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(19),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][19]~q\);

-- Location: LABCELL_X56_Y1_N12
\RegFile[10][19]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[10][19]~feeder_combout\ = ( \R.regWriteData\(19) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(19),
	combout => \RegFile[10][19]~feeder_combout\);

-- Location: FF_X56_Y1_N13
\RegFile[10][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[10][19]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][19]~q\);

-- Location: LABCELL_X63_Y1_N30
\RegFile[11][19]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[11][19]~feeder_combout\ = ( \R.regWriteData\(19) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(19),
	combout => \RegFile[11][19]~feeder_combout\);

-- Location: FF_X63_Y1_N32
\RegFile[11][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[11][19]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][19]~q\);

-- Location: FF_X66_Y5_N49
\RegFile[8][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(19),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][19]~q\);

-- Location: LABCELL_X63_Y1_N0
\Mux103~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux103~14_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[8][19]~q\))) # (\R.curInst\(20) & (\RegFile[9][19]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & (\RegFile[10][19]~q\)) # (\R.curInst\(20) & ((\RegFile[11][19]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][19]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[10][19]~q\,
	datad => \ALT_INV_RegFile[11][19]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][19]~q\,
	combout => \Mux103~14_combout\);

-- Location: FF_X63_Y3_N7
\RegFile[12][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(19),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][19]~q\);

-- Location: LABCELL_X63_Y1_N54
\Mux103~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux103~1_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux103~14_combout\)))) # (\R.curInst\(22) & ((!\Mux103~14_combout\ & ((\RegFile[12][19]~q\))) # (\Mux103~14_combout\ & (\RegFile[13][19]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux103~14_combout\)))) # (\R.curInst\(22) & ((!\Mux103~14_combout\ & ((\RegFile[14][19]~q\))) # (\Mux103~14_combout\ & (\RegFile[15][19]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][19]~q\,
	datab => \ALT_INV_RegFile[15][19]~q\,
	datac => \ALT_INV_RegFile[14][19]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux103~14_combout\,
	datag => \ALT_INV_RegFile[12][19]~q\,
	combout => \Mux103~1_combout\);

-- Location: LABCELL_X74_Y1_N12
\Mux103~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux103~13_combout\ = ( \Mux103~9_combout\ & ( \Mux103~1_combout\ & ( ((!\R.curInst\(24) & ((\Mux103~26_combout\))) # (\R.curInst\(24) & (\Mux103~5_combout\))) # (\R.curInst\(23)) ) ) ) # ( !\Mux103~9_combout\ & ( \Mux103~1_combout\ & ( (!\R.curInst\(23) 
-- & ((!\R.curInst\(24) & ((\Mux103~26_combout\))) # (\R.curInst\(24) & (\Mux103~5_combout\)))) # (\R.curInst\(23) & (!\R.curInst\(24))) ) ) ) # ( \Mux103~9_combout\ & ( !\Mux103~1_combout\ & ( (!\R.curInst\(23) & ((!\R.curInst\(24) & 
-- ((\Mux103~26_combout\))) # (\R.curInst\(24) & (\Mux103~5_combout\)))) # (\R.curInst\(23) & (\R.curInst\(24))) ) ) ) # ( !\Mux103~9_combout\ & ( !\Mux103~1_combout\ & ( (!\R.curInst\(23) & ((!\R.curInst\(24) & ((\Mux103~26_combout\))) # (\R.curInst\(24) & 
-- (\Mux103~5_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001010001010000100111001101101000110110011100101011111011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(23),
	datab => \ALT_INV_R.curInst\(24),
	datac => \ALT_INV_Mux103~5_combout\,
	datad => \ALT_INV_Mux103~26_combout\,
	datae => \ALT_INV_Mux103~9_combout\,
	dataf => \ALT_INV_Mux103~1_combout\,
	combout => \Mux103~13_combout\);

-- Location: LABCELL_X75_Y4_N15
\NxR.aluData2[19]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[19]~2_combout\ = ( \Mux103~13_combout\ & ( (!\vAluSrc2~1_combout\) # ((\Equal4~1_combout\ & \Mux135~0_combout\)) ) ) # ( !\Mux103~13_combout\ & ( (\Equal4~1_combout\ & (\vAluSrc2~1_combout\ & \Mux135~0_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000101000000000000010111110000111101011111000011110101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Equal4~1_combout\,
	datac => \ALT_INV_vAluSrc2~1_combout\,
	datad => \ALT_INV_Mux135~0_combout\,
	dataf => \ALT_INV_Mux103~13_combout\,
	combout => \NxR.aluData2[19]~2_combout\);

-- Location: FF_X75_Y4_N17
\R.aluData2[19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR.aluData2[19]~2_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData2\(19));

-- Location: LABCELL_X77_Y6_N0
\Selector13~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector13~4_combout\ = ( \R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( (!\R.aluData1\(19) & ((!\R.aluData2\(19)) # ((!\R.aluOp.ALUOpXor~DUPLICATE_q\ & !\R.aluOp.ALUOpOr~q\)))) # (\R.aluData1\(19) & (!\R.aluData2\(19) & (!\R.aluOp.ALUOpXor~DUPLICATE_q\ & 
-- !\R.aluOp.ALUOpOr~q\))) ) ) # ( !\R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( (!\R.aluOp.ALUOpOr~q\ & ((!\R.aluOp.ALUOpXor~DUPLICATE_q\) # (!\R.aluData1\(19) $ (\R.aluData2\(19))))) # (\R.aluOp.ALUOpOr~q\ & (!\R.aluData1\(19) & (!\R.aluData2\(19)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111100110001000111110011000100011101000100010001110100010001000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData1\(19),
	datab => \ALT_INV_R.aluData2\(19),
	datac => \ALT_INV_R.aluOp.ALUOpXor~DUPLICATE_q\,
	datad => \ALT_INV_R.aluOp.ALUOpOr~q\,
	dataf => \ALT_INV_R.aluOp.ALUOpAnd~DUPLICATE_q\,
	combout => \Selector13~4_combout\);

-- Location: LABCELL_X79_Y5_N57
\Selector13~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector13~5_combout\ = ( \Selector13~4_combout\ & ( (!\Selector16~0_OTERM393\) # (!\ShiftLeft0~3_OTERM223\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111100001111111111110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Selector16~0_OTERM393\,
	datad => \ALT_INV_ShiftLeft0~3_OTERM223\,
	dataf => \ALT_INV_Selector13~4_combout\,
	combout => \Selector13~5_combout\);

-- Location: LABCELL_X75_Y4_N42
\Mux136~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux136~0_combout\ = ( \Mux123~2_combout\ & ( \R.curInst\(18) ) ) # ( !\Mux123~2_combout\ & ( \R.curInst\(18) & ( ((\vAluSrc1~0_combout\ & ((\R.curInst\(2)) # (\Mux124~0_combout\)))) # (\Mux149~0_combout\) ) ) ) # ( \Mux123~2_combout\ & ( !\R.curInst\(18) 
-- ) ) # ( !\Mux123~2_combout\ & ( !\R.curInst\(18) & ( (\Mux124~0_combout\ & \vAluSrc1~0_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010101111111111111111100001111011111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux124~0_combout\,
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_Mux149~0_combout\,
	datad => \ALT_INV_vAluSrc1~0_combout\,
	datae => \ALT_INV_Mux123~2_combout\,
	dataf => \ALT_INV_R.curInst\(18),
	combout => \Mux136~0_combout\);

-- Location: FF_X65_Y5_N50
\RegFile[15][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(18),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][18]~q\);

-- Location: FF_X65_Y5_N32
\RegFile[13][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(18),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][18]~q\);

-- Location: MLABCELL_X65_Y5_N57
\RegFile[14][18]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[14][18]~feeder_combout\ = ( \R.regWriteData\(18) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(18),
	combout => \RegFile[14][18]~feeder_combout\);

-- Location: FF_X65_Y5_N58
\RegFile[14][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[14][18]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][18]~q\);

-- Location: FF_X65_Y3_N20
\RegFile[9][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(18),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][18]~q\);

-- Location: MLABCELL_X65_Y3_N54
\RegFile[10][18]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[10][18]~feeder_combout\ = ( \R.regWriteData\(18) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(18),
	combout => \RegFile[10][18]~feeder_combout\);

-- Location: FF_X65_Y3_N55
\RegFile[10][18]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[10][18]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][18]~DUPLICATE_q\);

-- Location: FF_X65_Y3_N26
\RegFile[11][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(18),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][18]~q\);

-- Location: LABCELL_X66_Y5_N39
\RegFile[8][18]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[8][18]~feeder_combout\ = ( \R.regWriteData\(18) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(18),
	combout => \RegFile[8][18]~feeder_combout\);

-- Location: FF_X66_Y5_N41
\RegFile[8][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[8][18]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][18]~q\);

-- Location: MLABCELL_X65_Y5_N42
\Mux104~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux104~14_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[8][18]~q\))) # (\R.curInst\(20) & (\RegFile[9][18]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & (\RegFile[10][18]~DUPLICATE_q\)) # (\R.curInst\(20) & ((\RegFile[11][18]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][18]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[10][18]~DUPLICATE_q\,
	datad => \ALT_INV_RegFile[11][18]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][18]~q\,
	combout => \Mux104~14_combout\);

-- Location: FF_X61_Y7_N40
\RegFile[12][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(18),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][18]~q\);

-- Location: MLABCELL_X65_Y5_N30
\Mux104~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux104~1_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux104~14_combout\)))) # (\R.curInst\(22) & ((!\Mux104~14_combout\ & ((\RegFile[12][18]~q\))) # (\Mux104~14_combout\ & (\RegFile[13][18]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux104~14_combout\)))) # (\R.curInst\(22) & ((!\Mux104~14_combout\ & ((\RegFile[14][18]~q\))) # (\Mux104~14_combout\ & (\RegFile[15][18]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][18]~q\,
	datab => \ALT_INV_RegFile[13][18]~q\,
	datac => \ALT_INV_RegFile[14][18]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux104~14_combout\,
	datag => \ALT_INV_RegFile[12][18]~q\,
	combout => \Mux104~1_combout\);

-- Location: FF_X64_Y4_N14
\RegFile[23][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(18),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][18]~q\);

-- Location: LABCELL_X64_Y4_N54
\RegFile[22][18]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[22][18]~feeder_combout\ = ( \R.regWriteData\(18) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(18),
	combout => \RegFile[22][18]~feeder_combout\);

-- Location: FF_X64_Y4_N55
\RegFile[22][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[22][18]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][18]~q\);

-- Location: FF_X64_Y4_N26
\RegFile[19][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(18),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][18]~q\);

-- Location: FF_X63_Y5_N4
\RegFile[18][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(18),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][18]~q\);

-- Location: FF_X63_Y5_N31
\RegFile[17][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(18),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][18]~q\);

-- Location: FF_X63_Y5_N47
\RegFile[16][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(18),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][18]~q\);

-- Location: MLABCELL_X65_Y7_N48
\Mux104~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux104~18_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & (\RegFile[16][18]~q\)) # (\R.curInst\(20) & ((\RegFile[17][18]~q\)))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & ((\RegFile[18][18]~q\))) # (\R.curInst\(20) & (\RegFile[19][18]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001010101111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[19][18]~q\,
	datac => \ALT_INV_RegFile[18][18]~q\,
	datad => \ALT_INV_RegFile[17][18]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][18]~q\,
	combout => \Mux104~18_combout\);

-- Location: LABCELL_X68_Y7_N18
\RegFile[20][18]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[20][18]~feeder_combout\ = ( \R.regWriteData\(18) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(18),
	combout => \RegFile[20][18]~feeder_combout\);

-- Location: FF_X68_Y7_N19
\RegFile[20][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[20][18]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][18]~q\);

-- Location: LABCELL_X68_Y7_N30
\Mux104~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux104~5_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux104~18_combout\)))) # (\R.curInst\(22) & ((!\Mux104~18_combout\ & (\RegFile[20][18]~q\)) # (\Mux104~18_combout\ & ((\RegFile[21][18]~q\)))))) ) ) # ( \R.curInst\(21) & ( 
-- (!\R.curInst\(22) & ((((\Mux104~18_combout\))))) # (\R.curInst\(22) & (((!\Mux104~18_combout\ & ((\RegFile[22][18]~q\))) # (\Mux104~18_combout\ & (\RegFile[23][18]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111001100111111111101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[23][18]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[22][18]~q\,
	datad => \ALT_INV_RegFile[21][18]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux104~18_combout\,
	datag => \ALT_INV_RegFile[20][18]~q\,
	combout => \Mux104~5_combout\);

-- Location: FF_X68_Y4_N8
\RegFile[3][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(18),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][18]~q\);

-- Location: FF_X68_Y7_N38
\RegFile[2][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(18),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][18]~q\);

-- Location: FF_X71_Y6_N44
\RegFile[5][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(18),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][18]~q\);

-- Location: FF_X67_Y5_N38
\RegFile[4][18]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(18),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][18]~DUPLICATE_q\);

-- Location: LABCELL_X68_Y4_N36
\RegFile[6][18]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[6][18]~feeder_combout\ = ( \R.regWriteData\(18) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(18),
	combout => \RegFile[6][18]~feeder_combout\);

-- Location: FF_X68_Y4_N37
\RegFile[6][18]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[6][18]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][18]~DUPLICATE_q\);

-- Location: FF_X68_Y4_N19
\RegFile[7][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(18),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][18]~q\);

-- Location: LABCELL_X68_Y7_N9
\Mux104~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux104~0_combout\ = ( \R.curInst\(20) & ( \R.curInst\(21) & ( \RegFile[7][18]~q\ ) ) ) # ( !\R.curInst\(20) & ( \R.curInst\(21) & ( \RegFile[6][18]~DUPLICATE_q\ ) ) ) # ( \R.curInst\(20) & ( !\R.curInst\(21) & ( \RegFile[5][18]~q\ ) ) ) # ( 
-- !\R.curInst\(20) & ( !\R.curInst\(21) & ( \RegFile[4][18]~DUPLICATE_q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110011010101010101010100001111000011110000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[5][18]~q\,
	datab => \ALT_INV_RegFile[4][18]~DUPLICATE_q\,
	datac => \ALT_INV_RegFile[6][18]~DUPLICATE_q\,
	datad => \ALT_INV_RegFile[7][18]~q\,
	datae => \ALT_INV_R.curInst\(20),
	dataf => \ALT_INV_R.curInst\(21),
	combout => \Mux104~0_combout\);

-- Location: LABCELL_X68_Y9_N24
\RegFile[1][18]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[1][18]~feeder_combout\ = ( \R.regWriteData\(18) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(18),
	combout => \RegFile[1][18]~feeder_combout\);

-- Location: FF_X68_Y9_N25
\RegFile[1][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[1][18]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][18]~q\);

-- Location: LABCELL_X68_Y7_N36
\Mux104~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux104~26_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (\RegFile[1][18]~q\ & (\R.curInst\(20)))) # (\R.curInst\(22) & (((\Mux104~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (((\RegFile[2][18]~q\)))) # 
-- (\R.curInst\(20) & (\RegFile[3][18]~q\)))) # (\R.curInst\(22) & ((((\Mux104~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001100000011000100010000110011001111110011111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][18]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[2][18]~q\,
	datad => \ALT_INV_R.curInst\(20),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux104~0_combout\,
	datag => \ALT_INV_RegFile[1][18]~q\,
	combout => \Mux104~26_combout\);

-- Location: FF_X62_Y6_N20
\RegFile[29][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(18),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][18]~q\);

-- Location: LABCELL_X62_Y6_N30
\RegFile[30][18]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[30][18]~feeder_combout\ = ( \R.regWriteData\(18) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(18),
	combout => \RegFile[30][18]~feeder_combout\);

-- Location: FF_X62_Y6_N31
\RegFile[30][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[30][18]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][18]~q\);

-- Location: FF_X62_Y4_N14
\RegFile[31][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(18),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][18]~q\);

-- Location: FF_X62_Y4_N8
\RegFile[25][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(18),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][18]~q\);

-- Location: LABCELL_X57_Y3_N48
\RegFile[26][18]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[26][18]~feeder_combout\ = ( \R.regWriteData\(18) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(18),
	combout => \RegFile[26][18]~feeder_combout\);

-- Location: FF_X57_Y3_N49
\RegFile[26][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[26][18]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][18]~q\);

-- Location: FF_X62_Y4_N50
\RegFile[27][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(18),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][18]~q\);

-- Location: LABCELL_X60_Y4_N24
\RegFile[24][18]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[24][18]~feeder_combout\ = ( \R.regWriteData\(18) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(18),
	combout => \RegFile[24][18]~feeder_combout\);

-- Location: FF_X60_Y4_N25
\RegFile[24][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[24][18]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][18]~q\);

-- Location: LABCELL_X62_Y4_N6
\Mux104~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux104~22_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[24][18]~q\))) # (\R.curInst\(20) & (\RegFile[25][18]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & (\RegFile[26][18]~q\)) # (\R.curInst\(20) & ((\RegFile[27][18]~q\)))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001110111011101110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[25][18]~q\,
	datac => \ALT_INV_RegFile[26][18]~q\,
	datad => \ALT_INV_RegFile[27][18]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][18]~q\,
	combout => \Mux104~22_combout\);

-- Location: LABCELL_X62_Y6_N12
\RegFile[28][18]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[28][18]~feeder_combout\ = ( \R.regWriteData\(18) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(18),
	combout => \RegFile[28][18]~feeder_combout\);

-- Location: FF_X62_Y6_N13
\RegFile[28][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[28][18]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][18]~q\);

-- Location: LABCELL_X62_Y6_N18
\Mux104~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux104~9_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux104~22_combout\))))) # (\R.curInst\(22) & (((!\Mux104~22_combout\ & ((\RegFile[28][18]~q\))) # (\Mux104~22_combout\ & (\RegFile[29][18]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux104~22_combout\)))) # (\R.curInst\(22) & ((!\Mux104~22_combout\ & (\RegFile[30][18]~q\)) # (\Mux104~22_combout\ & ((\RegFile[31][18]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[29][18]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[30][18]~q\,
	datad => \ALT_INV_RegFile[31][18]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux104~22_combout\,
	datag => \ALT_INV_RegFile[28][18]~q\,
	combout => \Mux104~9_combout\);

-- Location: LABCELL_X68_Y7_N24
\Mux104~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux104~13_combout\ = ( \Mux104~26_combout\ & ( \Mux104~9_combout\ & ( (!\R.curInst\(23) & (((!\R.curInst\(24)) # (\Mux104~5_combout\)))) # (\R.curInst\(23) & (((\R.curInst\(24))) # (\Mux104~1_combout\))) ) ) ) # ( !\Mux104~26_combout\ & ( 
-- \Mux104~9_combout\ & ( (!\R.curInst\(23) & (((\R.curInst\(24) & \Mux104~5_combout\)))) # (\R.curInst\(23) & (((\R.curInst\(24))) # (\Mux104~1_combout\))) ) ) ) # ( \Mux104~26_combout\ & ( !\Mux104~9_combout\ & ( (!\R.curInst\(23) & (((!\R.curInst\(24)) # 
-- (\Mux104~5_combout\)))) # (\R.curInst\(23) & (\Mux104~1_combout\ & (!\R.curInst\(24)))) ) ) ) # ( !\Mux104~26_combout\ & ( !\Mux104~9_combout\ & ( (!\R.curInst\(23) & (((\R.curInst\(24) & \Mux104~5_combout\)))) # (\R.curInst\(23) & (\Mux104~1_combout\ & 
-- (!\R.curInst\(24)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000000011010101100001011101000010101000111111011010110111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(23),
	datab => \ALT_INV_Mux104~1_combout\,
	datac => \ALT_INV_R.curInst\(24),
	datad => \ALT_INV_Mux104~5_combout\,
	datae => \ALT_INV_Mux104~26_combout\,
	dataf => \ALT_INV_Mux104~9_combout\,
	combout => \Mux104~13_combout\);

-- Location: LABCELL_X75_Y4_N33
\NxR.aluData2[18]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[18]~3_combout\ = ( \Mux104~13_combout\ & ( (!\vAluSrc2~1_combout\) # ((\Equal4~1_combout\ & \Mux136~0_combout\)) ) ) # ( !\Mux104~13_combout\ & ( (\Equal4~1_combout\ & (\vAluSrc2~1_combout\ & \Mux136~0_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000101000000000000010111110000111101011111000011110101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Equal4~1_combout\,
	datac => \ALT_INV_vAluSrc2~1_combout\,
	datad => \ALT_INV_Mux136~0_combout\,
	dataf => \ALT_INV_Mux104~13_combout\,
	combout => \NxR.aluData2[18]~3_combout\);

-- Location: FF_X75_Y4_N35
\R.aluData2[18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR.aluData2[18]~3_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData2\(18));

-- Location: FF_X74_Y6_N52
\Add2~65_OTERM703_NEW_REG804\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux237~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Add2~65_OTERM703_OTERM805\);

-- Location: LABCELL_X75_Y4_N54
\Mux138~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux138~0_combout\ = ( \Mux123~2_combout\ & ( \R.curInst\(16) ) ) # ( !\Mux123~2_combout\ & ( \R.curInst\(16) & ( ((\vAluSrc1~0_combout\ & ((\R.curInst\(2)) # (\Mux124~0_combout\)))) # (\Mux149~0_combout\) ) ) ) # ( \Mux123~2_combout\ & ( !\R.curInst\(16) 
-- ) ) # ( !\Mux123~2_combout\ & ( !\R.curInst\(16) & ( (\Mux124~0_combout\ & \vAluSrc1~0_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010101111111111111111100001111011111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux124~0_combout\,
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_Mux149~0_combout\,
	datad => \ALT_INV_vAluSrc1~0_combout\,
	datae => \ALT_INV_Mux123~2_combout\,
	dataf => \ALT_INV_R.curInst\(16),
	combout => \Mux138~0_combout\);

-- Location: LABCELL_X81_Y6_N42
\Add0~57\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~57_sumout\ = SUM(( \R.curPC\(16) ) + ( GND ) + ( \Add0~54\ ))
-- \Add0~58\ = CARRY(( \R.curPC\(16) ) + ( GND ) + ( \Add0~54\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.curPC\(16),
	cin => \Add0~54\,
	sumout => \Add0~57_sumout\,
	cout => \Add0~58\);

-- Location: LABCELL_X79_Y3_N51
\R.regWriteData[16]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.regWriteData[16]~feeder_combout\ = ( \Add0~57_sumout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_Add0~57_sumout\,
	combout => \R.regWriteData[16]~feeder_combout\);

-- Location: FF_X73_Y6_N10
\Add2~65_OTERM703_NEW_REG808\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux238~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Add2~65_OTERM703_OTERM809\);

-- Location: MLABCELL_X78_Y6_N42
\Add1~57\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~57_sumout\ = SUM(( \Add2~57_OTERM707_OTERM813\ ) + ( \Add2~57_OTERM707_OTERM815\ ) + ( \Add1~54\ ))
-- \Add1~58\ = CARRY(( \Add2~57_OTERM707_OTERM813\ ) + ( \Add2~57_OTERM707_OTERM815\ ) + ( \Add1~54\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Add2~57_OTERM707_OTERM815\,
	datad => \ALT_INV_Add2~57_OTERM707_OTERM813\,
	cin => \Add1~54\,
	sumout => \Add1~57_sumout\,
	cout => \Add1~58\);

-- Location: MLABCELL_X78_Y6_N45
\Add1~61\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~61_sumout\ = SUM(( \R.aluData1\(15) ) + ( \R.aluData2\(15) ) + ( \Add1~58\ ))
-- \Add1~62\ = CARRY(( \R.aluData1\(15) ) + ( \R.aluData2\(15) ) + ( \Add1~58\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluData2\(15),
	datad => \ALT_INV_R.aluData1\(15),
	cin => \Add1~58\,
	sumout => \Add1~61_sumout\,
	cout => \Add1~62\);

-- Location: MLABCELL_X78_Y6_N48
\Add1~65\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~65_sumout\ = SUM(( \Add2~65_OTERM703_OTERM811\ ) + ( \Add2~65_OTERM703_OTERM809\ ) + ( \Add1~62\ ))
-- \Add1~66\ = CARRY(( \Add2~65_OTERM703_OTERM811\ ) + ( \Add2~65_OTERM703_OTERM809\ ) + ( \Add1~62\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Add2~65_OTERM703_OTERM811\,
	datac => \ALT_INV_Add2~65_OTERM703_OTERM809\,
	cin => \Add1~62\,
	sumout => \Add1~65_sumout\,
	cout => \Add1~66\);

-- Location: FF_X73_Y7_N4
\Add2~25_OTERM723_NEW_REG832\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux248~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Add2~25_OTERM723_OTERM833\);

-- Location: LABCELL_X79_Y6_N18
\Add2~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~25_sumout\ = SUM(( !\Add2~25_OTERM723_OTERM835\ $ (\Add2~25_OTERM723_OTERM833\) ) + ( \Add2~23\ ) + ( \Add2~22\ ))
-- \Add2~26\ = CARRY(( !\Add2~25_OTERM723_OTERM835\ $ (\Add2~25_OTERM723_OTERM833\) ) + ( \Add2~23\ ) + ( \Add2~22\ ))
-- \Add2~27\ = SHARE((!\Add2~25_OTERM723_OTERM835\ & \Add2~25_OTERM723_OTERM833\))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000001111000000000000000000001111000000001111",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Add2~25_OTERM723_OTERM835\,
	datad => \ALT_INV_Add2~25_OTERM723_OTERM833\,
	cin => \Add2~22\,
	sharein => \Add2~23\,
	sumout => \Add2~25_sumout\,
	cout => \Add2~26\,
	shareout => \Add2~27\);

-- Location: LABCELL_X79_Y6_N21
\Add2~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~29_sumout\ = SUM(( !\Add2~25_OTERM723_OTERM829\ $ (\Add2~25_OTERM723_OTERM831\) ) + ( \Add2~27\ ) + ( \Add2~26\ ))
-- \Add2~30\ = CARRY(( !\Add2~25_OTERM723_OTERM829\ $ (\Add2~25_OTERM723_OTERM831\) ) + ( \Add2~27\ ) + ( \Add2~26\ ))
-- \Add2~31\ = SHARE((\Add2~25_OTERM723_OTERM829\ & !\Add2~25_OTERM723_OTERM831\))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000000000000000000000001111000000001111",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Add2~25_OTERM723_OTERM829\,
	datad => \ALT_INV_Add2~25_OTERM723_OTERM831\,
	cin => \Add2~26\,
	sharein => \Add2~27\,
	sumout => \Add2~29_sumout\,
	cout => \Add2~30\,
	shareout => \Add2~31\);

-- Location: LABCELL_X79_Y6_N24
\Add2~33\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~33_sumout\ = SUM(( !\Add2~33_OTERM719_OTERM827\ $ (\Add2~33_OTERM719_OTERM825\) ) + ( \Add2~31\ ) + ( \Add2~30\ ))
-- \Add2~34\ = CARRY(( !\Add2~33_OTERM719_OTERM827\ $ (\Add2~33_OTERM719_OTERM825\) ) + ( \Add2~31\ ) + ( \Add2~30\ ))
-- \Add2~35\ = SHARE((!\Add2~33_OTERM719_OTERM827\ & \Add2~33_OTERM719_OTERM825\))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000001111000000000000000000001111000000001111",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Add2~33_OTERM719_OTERM827\,
	datad => \ALT_INV_Add2~33_OTERM719_OTERM825\,
	cin => \Add2~30\,
	sharein => \Add2~31\,
	sumout => \Add2~33_sumout\,
	cout => \Add2~34\,
	shareout => \Add2~35\);

-- Location: LABCELL_X79_Y6_N27
\Add2~37\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~37_sumout\ = SUM(( !\Add2~33_OTERM719_OTERM823\ $ (\Add2~33_OTERM719_OTERM821\) ) + ( \Add2~35\ ) + ( \Add2~34\ ))
-- \Add2~38\ = CARRY(( !\Add2~33_OTERM719_OTERM823\ $ (\Add2~33_OTERM719_OTERM821\) ) + ( \Add2~35\ ) + ( \Add2~34\ ))
-- \Add2~39\ = SHARE((!\Add2~33_OTERM719_OTERM823\ & \Add2~33_OTERM719_OTERM821\))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011000000110000000000000000001100001111000011",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Add2~33_OTERM719_OTERM823\,
	datac => \ALT_INV_Add2~33_OTERM719_OTERM821\,
	cin => \Add2~34\,
	sharein => \Add2~35\,
	sumout => \Add2~37_sumout\,
	cout => \Add2~38\,
	shareout => \Add2~39\);

-- Location: LABCELL_X79_Y6_N30
\Add2~41\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~41_sumout\ = SUM(( !\Add2~41_OTERM715_OTERM819\ $ (\Add2~41_OTERM715_OTERM817\) ) + ( \Add2~39\ ) + ( \Add2~38\ ))
-- \Add2~42\ = CARRY(( !\Add2~41_OTERM715_OTERM819\ $ (\Add2~41_OTERM715_OTERM817\) ) + ( \Add2~39\ ) + ( \Add2~38\ ))
-- \Add2~43\ = SHARE((!\Add2~41_OTERM715_OTERM819\ & \Add2~41_OTERM715_OTERM817\))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000001111000000000000000000001111000000001111",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Add2~41_OTERM715_OTERM819\,
	datad => \ALT_INV_Add2~41_OTERM715_OTERM817\,
	cin => \Add2~38\,
	sharein => \Add2~39\,
	sumout => \Add2~41_sumout\,
	cout => \Add2~42\,
	shareout => \Add2~43\);

-- Location: LABCELL_X79_Y6_N33
\Add2~45\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~45_sumout\ = SUM(( !\R.aluData2\(11) $ (\R.aluData1\(11)) ) + ( \Add2~43\ ) + ( \Add2~42\ ))
-- \Add2~46\ = CARRY(( !\R.aluData2\(11) $ (\R.aluData1\(11)) ) + ( \Add2~43\ ) + ( \Add2~42\ ))
-- \Add2~47\ = SHARE((!\R.aluData2\(11) & \R.aluData1\(11)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000001010101000000000000000001010101001010101",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(11),
	datad => \ALT_INV_R.aluData1\(11),
	cin => \Add2~42\,
	sharein => \Add2~43\,
	sumout => \Add2~45_sumout\,
	cout => \Add2~46\,
	shareout => \Add2~47\);

-- Location: LABCELL_X79_Y6_N36
\Add2~49\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~49_sumout\ = SUM(( !\R.aluData1\(12) $ (\R.aluData2\(12)) ) + ( \Add2~47\ ) + ( \Add2~46\ ))
-- \Add2~50\ = CARRY(( !\R.aluData1\(12) $ (\R.aluData2\(12)) ) + ( \Add2~47\ ) + ( \Add2~46\ ))
-- \Add2~51\ = SHARE((\R.aluData1\(12) & !\R.aluData2\(12)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000000000000000000000001111000000001111",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluData1\(12),
	datad => \ALT_INV_R.aluData2\(12),
	cin => \Add2~46\,
	sharein => \Add2~47\,
	sumout => \Add2~49_sumout\,
	cout => \Add2~50\,
	shareout => \Add2~51\);

-- Location: LABCELL_X79_Y6_N39
\Add2~53\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~53_sumout\ = SUM(( !\R.aluData2\(13) $ (\R.aluData1\(13)) ) + ( \Add2~51\ ) + ( \Add2~50\ ))
-- \Add2~54\ = CARRY(( !\R.aluData2\(13) $ (\R.aluData1\(13)) ) + ( \Add2~51\ ) + ( \Add2~50\ ))
-- \Add2~55\ = SHARE((!\R.aluData2\(13) & \R.aluData1\(13)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000001111000000000000000000001111000000001111",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluData2\(13),
	datad => \ALT_INV_R.aluData1\(13),
	cin => \Add2~50\,
	sharein => \Add2~51\,
	sumout => \Add2~53_sumout\,
	cout => \Add2~54\,
	shareout => \Add2~55\);

-- Location: LABCELL_X79_Y6_N42
\Add2~57\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~57_sumout\ = SUM(( !\Add2~57_OTERM707_OTERM815\ $ (\Add2~57_OTERM707_OTERM813\) ) + ( \Add2~55\ ) + ( \Add2~54\ ))
-- \Add2~58\ = CARRY(( !\Add2~57_OTERM707_OTERM815\ $ (\Add2~57_OTERM707_OTERM813\) ) + ( \Add2~55\ ) + ( \Add2~54\ ))
-- \Add2~59\ = SHARE((!\Add2~57_OTERM707_OTERM815\ & \Add2~57_OTERM707_OTERM813\))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011000000110000000000000000001100001111000011",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Add2~57_OTERM707_OTERM815\,
	datac => \ALT_INV_Add2~57_OTERM707_OTERM813\,
	cin => \Add2~54\,
	sharein => \Add2~55\,
	sumout => \Add2~57_sumout\,
	cout => \Add2~58\,
	shareout => \Add2~59\);

-- Location: LABCELL_X79_Y6_N45
\Add2~61\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~61_sumout\ = SUM(( !\R.aluData2\(15) $ (\R.aluData1\(15)) ) + ( \Add2~59\ ) + ( \Add2~58\ ))
-- \Add2~62\ = CARRY(( !\R.aluData2\(15) $ (\R.aluData1\(15)) ) + ( \Add2~59\ ) + ( \Add2~58\ ))
-- \Add2~63\ = SHARE((!\R.aluData2\(15) & \R.aluData1\(15)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000001010101000000000000000001010101001010101",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(15),
	datad => \ALT_INV_R.aluData1\(15),
	cin => \Add2~58\,
	sharein => \Add2~59\,
	sumout => \Add2~61_sumout\,
	cout => \Add2~62\,
	shareout => \Add2~63\);

-- Location: LABCELL_X79_Y6_N48
\Add2~65\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~65_sumout\ = SUM(( !\Add2~65_OTERM703_OTERM809\ $ (\Add2~65_OTERM703_OTERM811\) ) + ( \Add2~63\ ) + ( \Add2~62\ ))
-- \Add2~66\ = CARRY(( !\Add2~65_OTERM703_OTERM809\ $ (\Add2~65_OTERM703_OTERM811\) ) + ( \Add2~63\ ) + ( \Add2~62\ ))
-- \Add2~67\ = SHARE((\Add2~65_OTERM703_OTERM809\ & !\Add2~65_OTERM703_OTERM811\))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000001100000011000000000000000000001100001111000011",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Add2~65_OTERM703_OTERM809\,
	datac => \ALT_INV_Add2~65_OTERM703_OTERM811\,
	cin => \Add2~62\,
	sharein => \Add2~63\,
	sumout => \Add2~65_sumout\,
	cout => \Add2~66\,
	shareout => \Add2~67\);

-- Location: LABCELL_X79_Y1_N21
\Comb:vRegWriteData[24]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[24]~1_combout\ = ( !\R.curInst\(14) & ( \R.memToReg~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.memToReg~q\,
	dataf => \ALT_INV_R.curInst\(14),
	combout => \Comb:vRegWriteData[24]~1_combout\);

-- Location: FF_X82_Y4_N2
\R.aluRes[16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector16~5_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(16));

-- Location: IOIBUF_X84_Y0_N18
\avm_d_readdata[23]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(23),
	o => \avm_d_readdata[23]~input_o\);

-- Location: IOIBUF_X84_Y0_N35
\avm_d_readdata[31]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(31),
	o => \avm_d_readdata[31]~input_o\);

-- Location: IOIBUF_X60_Y0_N1
\avm_d_readdata[8]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(8),
	o => \avm_d_readdata[8]~input_o\);

-- Location: LABCELL_X79_Y2_N18
\Comb:vRegWriteData[16]~0_RESYN1724\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[16]~0_RESYN1724_BDD1725\ = ( \R.curInst\(12) & ( (\avm_d_readdata[23]~input_o\ & !\R.curInst\(13)) ) ) # ( !\R.curInst\(12) & ( (!\R.curInst\(13) & (\avm_d_readdata[31]~input_o\)) # (\R.curInst\(13) & ((\avm_d_readdata[8]~input_o\))) ) 
-- )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011000000111111001100000011111101010000010100000101000001010000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_avm_d_readdata[23]~input_o\,
	datab => \ALT_INV_avm_d_readdata[31]~input_o\,
	datac => \ALT_INV_R.curInst\(13),
	datad => \ALT_INV_avm_d_readdata[8]~input_o\,
	dataf => \ALT_INV_R.curInst\(12),
	combout => \Comb:vRegWriteData[16]~0_RESYN1724_BDD1725\);

-- Location: LABCELL_X79_Y3_N48
\Comb:vRegWriteData[16]~0_RESYN1726\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[16]~0_RESYN1726_BDD1727\ = ( \Comb:vRegWriteData[16]~0_RESYN1724_BDD1725\ & ( ((!\R.aluCalc~q\ & (\R.aluRes\(16) & !\R.memToReg~q\))) # (\Comb:vRegWriteData[24]~1_combout\) ) ) # ( !\Comb:vRegWriteData[16]~0_RESYN1724_BDD1725\ & ( 
-- (!\R.aluCalc~q\ & (\R.aluRes\(16) & !\R.memToReg~q\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000110000000000000011000000000001011101010101010101110101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Comb:vRegWriteData[24]~1_combout\,
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_R.aluRes\(16),
	datad => \ALT_INV_R.memToReg~q\,
	dataf => \ALT_INV_Comb:vRegWriteData[16]~0_RESYN1724_BDD1725\,
	combout => \Comb:vRegWriteData[16]~0_RESYN1726_BDD1727\);

-- Location: LABCELL_X79_Y3_N15
\Comb:vRegWriteData[16]~0_RESYN1728\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[16]~0_RESYN1728_BDD1729\ = ( \R.memToReg~q\ & ( \Comb:vRegWriteData[16]~0_RESYN1726_BDD1727\ ) ) # ( !\R.memToReg~q\ & ( \Comb:vRegWriteData[16]~0_RESYN1726_BDD1727\ ) ) # ( !\R.memToReg~q\ & ( 
-- !\Comb:vRegWriteData[16]~0_RESYN1726_BDD1727\ & ( (\R.aluOp.ALUOpSub~q\ & (\Add2~65_sumout\ & \R.aluCalc~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000011000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_Add2~65_sumout\,
	datad => \ALT_INV_R.aluCalc~q\,
	datae => \ALT_INV_R.memToReg~q\,
	dataf => \ALT_INV_Comb:vRegWriteData[16]~0_RESYN1726_BDD1727\,
	combout => \Comb:vRegWriteData[16]~0_RESYN1728_BDD1729\);

-- Location: LABCELL_X79_Y3_N54
\Comb:vRegWriteData[16]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[16]~0_combout\ = ( \Add1~65_sumout\ & ( \Comb:vRegWriteData[16]~0_RESYN1728_BDD1729\ ) ) # ( !\Add1~65_sumout\ & ( \Comb:vRegWriteData[16]~0_RESYN1728_BDD1729\ ) ) # ( \Add1~65_sumout\ & ( !\Comb:vRegWriteData[16]~0_RESYN1728_BDD1729\ 
-- & ( (\R.aluCalc~q\ & (!\R.memToReg~q\ & ((!\Selector16~3_combout\) # (\R.aluOp.ALUOpAdd~q\)))) ) ) ) # ( !\Add1~65_sumout\ & ( !\Comb:vRegWriteData[16]~0_RESYN1728_BDD1729\ & ( (\R.aluCalc~q\ & (!\Selector16~3_combout\ & !\R.memToReg~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100010000000000010001010000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluCalc~q\,
	datab => \ALT_INV_Selector16~3_combout\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_R.memToReg~q\,
	datae => \ALT_INV_Add1~65_sumout\,
	dataf => \ALT_INV_Comb:vRegWriteData[16]~0_RESYN1728_BDD1729\,
	combout => \Comb:vRegWriteData[16]~0_combout\);

-- Location: FF_X79_Y3_N53
\R.regWriteData[16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \R.regWriteData[16]~feeder_combout\,
	asdata => \Comb:vRegWriteData[16]~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(16));

-- Location: FF_X65_Y2_N56
\RegFile[23][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][16]~q\);

-- Location: FF_X71_Y1_N14
\RegFile[21][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][16]~q\);

-- Location: FF_X71_Y1_N8
\RegFile[22][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][16]~q\);

-- Location: FF_X65_Y2_N20
\RegFile[19][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][16]~q\);

-- Location: FF_X63_Y5_N10
\RegFile[18][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][16]~q\);

-- Location: FF_X65_Y2_N32
\RegFile[17][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][16]~q\);

-- Location: FF_X63_Y5_N43
\RegFile[16][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][16]~q\);

-- Location: MLABCELL_X65_Y2_N30
\Mux106~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux106~18_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & (\RegFile[16][16]~q\)) # (\R.curInst\(20) & ((\RegFile[17][16]~q\)))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & ((\RegFile[18][16]~q\))) # (\R.curInst\(20) & (\RegFile[19][16]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001010101111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[19][16]~q\,
	datac => \ALT_INV_RegFile[18][16]~q\,
	datad => \ALT_INV_RegFile[17][16]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][16]~q\,
	combout => \Mux106~18_combout\);

-- Location: FF_X71_Y1_N56
\RegFile[20][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][16]~q\);

-- Location: LABCELL_X71_Y1_N42
\Mux106~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux106~5_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux106~18_combout\)))) # (\R.curInst\(22) & ((!\Mux106~18_combout\ & ((\RegFile[20][16]~q\))) # (\Mux106~18_combout\ & (\RegFile[21][16]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux106~18_combout\)))) # (\R.curInst\(22) & ((!\Mux106~18_combout\ & ((\RegFile[22][16]~q\))) # (\Mux106~18_combout\ & (\RegFile[23][16]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[23][16]~q\,
	datab => \ALT_INV_RegFile[21][16]~q\,
	datac => \ALT_INV_RegFile[22][16]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux106~18_combout\,
	datag => \ALT_INV_RegFile[20][16]~q\,
	combout => \Mux106~5_combout\);

-- Location: FF_X63_Y3_N14
\RegFile[15][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][16]~q\);

-- Location: FF_X63_Y3_N1
\RegFile[14][16]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][16]~DUPLICATE_q\);

-- Location: FF_X63_Y1_N50
\RegFile[13][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][16]~q\);

-- Location: FF_X63_Y1_N44
\RegFile[9][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][16]~q\);

-- Location: LABCELL_X60_Y2_N3
\RegFile[10][16]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[10][16]~feeder_combout\ = ( \R.regWriteData\(16) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(16),
	combout => \RegFile[10][16]~feeder_combout\);

-- Location: FF_X60_Y2_N4
\RegFile[10][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[10][16]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][16]~q\);

-- Location: FF_X63_Y1_N14
\RegFile[11][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][16]~q\);

-- Location: MLABCELL_X59_Y1_N42
\RegFile[8][16]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[8][16]~feeder_combout\ = ( \R.regWriteData\(16) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(16),
	combout => \RegFile[8][16]~feeder_combout\);

-- Location: FF_X59_Y1_N43
\RegFile[8][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[8][16]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][16]~q\);

-- Location: LABCELL_X63_Y1_N42
\Mux106~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux106~14_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[8][16]~q\))) # (\R.curInst\(20) & (\RegFile[9][16]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & (\RegFile[10][16]~q\)) # (\R.curInst\(20) & ((\RegFile[11][16]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][16]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[10][16]~q\,
	datad => \ALT_INV_RegFile[11][16]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][16]~q\,
	combout => \Mux106~14_combout\);

-- Location: FF_X63_Y3_N22
\RegFile[12][16]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][16]~DUPLICATE_q\);

-- Location: LABCELL_X63_Y1_N48
\Mux106~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux106~1_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux106~14_combout\)))) # (\R.curInst\(22) & ((!\Mux106~14_combout\ & (\RegFile[12][16]~DUPLICATE_q\)) # (\Mux106~14_combout\ & ((\RegFile[13][16]~q\)))))) ) ) # ( \R.curInst\(21) & ( 
-- (!\R.curInst\(22) & ((((\Mux106~14_combout\))))) # (\R.curInst\(22) & (((!\Mux106~14_combout\ & ((\RegFile[14][16]~DUPLICATE_q\))) # (\Mux106~14_combout\ & (\RegFile[15][16]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111001100111111111101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][16]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[14][16]~DUPLICATE_q\,
	datad => \ALT_INV_RegFile[13][16]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux106~14_combout\,
	datag => \ALT_INV_RegFile[12][16]~DUPLICATE_q\,
	combout => \Mux106~1_combout\);

-- Location: FF_X68_Y3_N44
\RegFile[3][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][16]~q\);

-- Location: FF_X72_Y3_N43
\RegFile[2][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][16]~q\);

-- Location: LABCELL_X67_Y5_N42
\RegFile[4][16]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[4][16]~feeder_combout\ = ( \R.regWriteData\(16) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(16),
	combout => \RegFile[4][16]~feeder_combout\);

-- Location: FF_X67_Y5_N43
\RegFile[4][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[4][16]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][16]~q\);

-- Location: FF_X68_Y3_N10
\RegFile[5][16]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][16]~DUPLICATE_q\);

-- Location: FF_X68_Y3_N49
\RegFile[7][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][16]~q\);

-- Location: FF_X71_Y3_N43
\RegFile[6][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][16]~q\);

-- Location: LABCELL_X71_Y3_N42
\Mux106~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux106~0_combout\ = ( \RegFile[6][16]~q\ & ( \R.curInst\(20) & ( (!\R.curInst\(21) & (\RegFile[5][16]~DUPLICATE_q\)) # (\R.curInst\(21) & ((\RegFile[7][16]~q\))) ) ) ) # ( !\RegFile[6][16]~q\ & ( \R.curInst\(20) & ( (!\R.curInst\(21) & 
-- (\RegFile[5][16]~DUPLICATE_q\)) # (\R.curInst\(21) & ((\RegFile[7][16]~q\))) ) ) ) # ( \RegFile[6][16]~q\ & ( !\R.curInst\(20) & ( (\R.curInst\(21)) # (\RegFile[4][16]~q\) ) ) ) # ( !\RegFile[6][16]~q\ & ( !\R.curInst\(20) & ( (\RegFile[4][16]~q\ & 
-- !\R.curInst\(21)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010100000000010101011111111100110011000011110011001100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[4][16]~q\,
	datab => \ALT_INV_RegFile[5][16]~DUPLICATE_q\,
	datac => \ALT_INV_RegFile[7][16]~q\,
	datad => \ALT_INV_R.curInst\(21),
	datae => \ALT_INV_RegFile[6][16]~q\,
	dataf => \ALT_INV_R.curInst\(20),
	combout => \Mux106~0_combout\);

-- Location: FF_X72_Y3_N38
\RegFile[1][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][16]~q\);

-- Location: LABCELL_X71_Y3_N12
\Mux106~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux106~26_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((\RegFile[1][16]~q\ & (\R.curInst\(20)))))) # (\R.curInst\(22) & ((((\Mux106~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (((\RegFile[2][16]~q\)))) 
-- # (\R.curInst\(20) & (\RegFile[3][16]~q\)))) # (\R.curInst\(22) & ((((\Mux106~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001010000010100010001001010101010111110101111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[3][16]~q\,
	datac => \ALT_INV_RegFile[2][16]~q\,
	datad => \ALT_INV_R.curInst\(20),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux106~0_combout\,
	datag => \ALT_INV_RegFile[1][16]~q\,
	combout => \Mux106~26_combout\);

-- Location: FF_X67_Y5_N2
\RegFile[31][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][16]~q\);

-- Location: LABCELL_X66_Y3_N36
\RegFile[30][16]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[30][16]~feeder_combout\ = \R.regWriteData\(16)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.regWriteData\(16),
	combout => \RegFile[30][16]~feeder_combout\);

-- Location: FF_X66_Y3_N37
\RegFile[30][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[30][16]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][16]~q\);

-- Location: FF_X66_Y2_N50
\RegFile[29][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][16]~q\);

-- Location: FF_X66_Y2_N26
\RegFile[25][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][16]~q\);

-- Location: LABCELL_X60_Y2_N42
\RegFile[26][16]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[26][16]~feeder_combout\ = ( \R.regWriteData\(16) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(16),
	combout => \RegFile[26][16]~feeder_combout\);

-- Location: FF_X60_Y2_N43
\RegFile[26][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[26][16]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][16]~q\);

-- Location: FF_X66_Y2_N14
\RegFile[27][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][16]~q\);

-- Location: MLABCELL_X59_Y2_N33
\RegFile[24][16]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[24][16]~feeder_combout\ = ( \R.regWriteData\(16) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(16),
	combout => \RegFile[24][16]~feeder_combout\);

-- Location: FF_X59_Y2_N34
\RegFile[24][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[24][16]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][16]~q\);

-- Location: LABCELL_X66_Y2_N24
\Mux106~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux106~22_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[24][16]~q\))) # (\R.curInst\(20) & (\RegFile[25][16]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & (\RegFile[26][16]~q\)) # (\R.curInst\(20) & ((\RegFile[27][16]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[25][16]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[26][16]~q\,
	datad => \ALT_INV_RegFile[27][16]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][16]~q\,
	combout => \Mux106~22_combout\);

-- Location: LABCELL_X66_Y3_N21
\RegFile[28][16]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[28][16]~feeder_combout\ = \R.regWriteData\(16)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101010101010101010101010101010101010101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.regWriteData\(16),
	combout => \RegFile[28][16]~feeder_combout\);

-- Location: FF_X66_Y3_N23
\RegFile[28][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[28][16]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][16]~q\);

-- Location: LABCELL_X66_Y2_N48
\Mux106~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux106~9_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux106~22_combout\))))) # (\R.curInst\(22) & (((!\Mux106~22_combout\ & (\RegFile[28][16]~q\)) # (\Mux106~22_combout\ & ((\RegFile[29][16]~q\)))))) ) ) # ( \R.curInst\(21) & ( 
-- (!\R.curInst\(22) & ((((\Mux106~22_combout\))))) # (\R.curInst\(22) & (((!\Mux106~22_combout\ & ((\RegFile[30][16]~q\))) # (\Mux106~22_combout\ & (\RegFile[31][16]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110101010111111111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[31][16]~q\,
	datac => \ALT_INV_RegFile[30][16]~q\,
	datad => \ALT_INV_RegFile[29][16]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux106~22_combout\,
	datag => \ALT_INV_RegFile[28][16]~q\,
	combout => \Mux106~9_combout\);

-- Location: LABCELL_X71_Y1_N33
\Mux106~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux106~13_combout\ = ( \Mux106~26_combout\ & ( \Mux106~9_combout\ & ( (!\R.curInst\(23) & (((!\R.curInst\(24))) # (\Mux106~5_combout\))) # (\R.curInst\(23) & (((\R.curInst\(24)) # (\Mux106~1_combout\)))) ) ) ) # ( !\Mux106~26_combout\ & ( 
-- \Mux106~9_combout\ & ( (!\R.curInst\(23) & (\Mux106~5_combout\ & ((\R.curInst\(24))))) # (\R.curInst\(23) & (((\R.curInst\(24)) # (\Mux106~1_combout\)))) ) ) ) # ( \Mux106~26_combout\ & ( !\Mux106~9_combout\ & ( (!\R.curInst\(23) & (((!\R.curInst\(24))) # 
-- (\Mux106~5_combout\))) # (\R.curInst\(23) & (((\Mux106~1_combout\ & !\R.curInst\(24))))) ) ) ) # ( !\Mux106~26_combout\ & ( !\Mux106~9_combout\ & ( (!\R.curInst\(23) & (\Mux106~5_combout\ & ((\R.curInst\(24))))) # (\R.curInst\(23) & (((\Mux106~1_combout\ 
-- & !\R.curInst\(24))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100100010101011110010001000000101011101111010111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(23),
	datab => \ALT_INV_Mux106~5_combout\,
	datac => \ALT_INV_Mux106~1_combout\,
	datad => \ALT_INV_R.curInst\(24),
	datae => \ALT_INV_Mux106~26_combout\,
	dataf => \ALT_INV_Mux106~9_combout\,
	combout => \Mux106~13_combout\);

-- Location: MLABCELL_X72_Y5_N48
\NxR.aluData2[16]~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[16]~5_combout\ = ( \Mux106~13_combout\ & ( (!\vAluSrc2~1_combout\) # ((\Equal4~1_combout\ & \Mux138~0_combout\)) ) ) # ( !\Mux106~13_combout\ & ( (\vAluSrc2~1_combout\ & (\Equal4~1_combout\ & \Mux138~0_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000010001000000000001000110101010101110111010101010111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluSrc2~1_combout\,
	datab => \ALT_INV_Equal4~1_combout\,
	datad => \ALT_INV_Mux138~0_combout\,
	dataf => \ALT_INV_Mux106~13_combout\,
	combout => \NxR.aluData2[16]~5_combout\);

-- Location: FF_X72_Y5_N59
\Add2~65_OTERM703_NEW_REG810\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \NxR.aluData2[16]~5_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Add2~65_OTERM703_OTERM811\);

-- Location: MLABCELL_X78_Y6_N51
\Add1~69\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~69_sumout\ = SUM(( \Add2~65_OTERM703_OTERM805\ ) + ( \Add2~65_OTERM703_OTERM807\ ) + ( \Add1~66\ ))
-- \Add1~70\ = CARRY(( \Add2~65_OTERM703_OTERM805\ ) + ( \Add2~65_OTERM703_OTERM807\ ) + ( \Add1~66\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Add2~65_OTERM703_OTERM807\,
	datad => \ALT_INV_Add2~65_OTERM703_OTERM805\,
	cin => \Add1~66\,
	sumout => \Add1~69_sumout\,
	cout => \Add1~70\);

-- Location: MLABCELL_X78_Y6_N54
\Add1~73\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~73_sumout\ = SUM(( \R.aluData1\(18) ) + ( \R.aluData2\(18) ) + ( \Add1~70\ ))
-- \Add1~74\ = CARRY(( \R.aluData1\(18) ) + ( \R.aluData2\(18) ) + ( \Add1~70\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluData2\(18),
	datad => \ALT_INV_R.aluData1\(18),
	cin => \Add1~70\,
	sumout => \Add1~73_sumout\,
	cout => \Add1~74\);

-- Location: MLABCELL_X78_Y6_N57
\Add1~77\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~77_sumout\ = SUM(( \R.aluData2\(19) ) + ( \R.aluData1\(19) ) + ( \Add1~74\ ))
-- \Add1~78\ = CARRY(( \R.aluData2\(19) ) + ( \R.aluData1\(19) ) + ( \Add1~74\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluData2\(19),
	dataf => \ALT_INV_R.aluData1\(19),
	cin => \Add1~74\,
	sumout => \Add1~77_sumout\,
	cout => \Add1~78\);

-- Location: LABCELL_X79_Y6_N51
\Add2~69\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~69_sumout\ = SUM(( !\Add2~65_OTERM703_OTERM807\ $ (\Add2~65_OTERM703_OTERM805\) ) + ( \Add2~67\ ) + ( \Add2~66\ ))
-- \Add2~70\ = CARRY(( !\Add2~65_OTERM703_OTERM807\ $ (\Add2~65_OTERM703_OTERM805\) ) + ( \Add2~67\ ) + ( \Add2~66\ ))
-- \Add2~71\ = SHARE((!\Add2~65_OTERM703_OTERM807\ & \Add2~65_OTERM703_OTERM805\))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000001111000000000000000000001111000000001111",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Add2~65_OTERM703_OTERM807\,
	datad => \ALT_INV_Add2~65_OTERM703_OTERM805\,
	cin => \Add2~66\,
	sharein => \Add2~67\,
	sumout => \Add2~69_sumout\,
	cout => \Add2~70\,
	shareout => \Add2~71\);

-- Location: LABCELL_X79_Y6_N54
\Add2~73\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~73_sumout\ = SUM(( !\R.aluData1\(18) $ (\R.aluData2\(18)) ) + ( \Add2~71\ ) + ( \Add2~70\ ))
-- \Add2~74\ = CARRY(( !\R.aluData1\(18) $ (\R.aluData2\(18)) ) + ( \Add2~71\ ) + ( \Add2~70\ ))
-- \Add2~75\ = SHARE((\R.aluData1\(18) & !\R.aluData2\(18)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000000000000000000000001111000000001111",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluData1\(18),
	datad => \ALT_INV_R.aluData2\(18),
	cin => \Add2~70\,
	sharein => \Add2~71\,
	sumout => \Add2~73_sumout\,
	cout => \Add2~74\,
	shareout => \Add2~75\);

-- Location: LABCELL_X79_Y6_N57
\Add2~77\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~77_sumout\ = SUM(( !\R.aluData1\(19) $ (\R.aluData2\(19)) ) + ( \Add2~75\ ) + ( \Add2~74\ ))
-- \Add2~78\ = CARRY(( !\R.aluData1\(19) $ (\R.aluData2\(19)) ) + ( \Add2~75\ ) + ( \Add2~74\ ))
-- \Add2~79\ = SHARE((\R.aluData1\(19) & !\R.aluData2\(19)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010101010000000000000000000000001010101001010101",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData1\(19),
	datad => \ALT_INV_R.aluData2\(19),
	cin => \Add2~74\,
	sharein => \Add2~75\,
	sumout => \Add2~77_sumout\,
	cout => \Add2~78\,
	shareout => \Add2~79\);

-- Location: LABCELL_X83_Y4_N18
\Selector13~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector13~1_combout\ = ( \Add1~77_sumout\ & ( \Add2~77_sumout\ & ( (\Selector13~5_combout\ & (!\R.aluOp.ALUOpSub~q\ & (!\R.aluOp.ALUOpAdd~q\ & !\Selector17~0_OTERM391\))) ) ) ) # ( !\Add1~77_sumout\ & ( \Add2~77_sumout\ & ( (\Selector13~5_combout\ & 
-- (!\R.aluOp.ALUOpSub~q\ & !\Selector17~0_OTERM391\)) ) ) ) # ( \Add1~77_sumout\ & ( !\Add2~77_sumout\ & ( (\Selector13~5_combout\ & (!\R.aluOp.ALUOpAdd~q\ & !\Selector17~0_OTERM391\)) ) ) ) # ( !\Add1~77_sumout\ & ( !\Add2~77_sumout\ & ( 
-- (\Selector13~5_combout\ & !\Selector17~0_OTERM391\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010100000000010100000000000001000100000000000100000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector13~5_combout\,
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_Selector17~0_OTERM391\,
	datae => \ALT_INV_Add1~77_sumout\,
	dataf => \ALT_INV_Add2~77_sumout\,
	combout => \Selector13~1_combout\);

-- Location: LABCELL_X79_Y5_N0
\Add2~81\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~81_sumout\ = SUM(( !\R.aluData2\(20) $ (\R.aluData1\(20)) ) + ( \Add2~79\ ) + ( \Add2~78\ ))
-- \Add2~82\ = CARRY(( !\R.aluData2\(20) $ (\R.aluData1\(20)) ) + ( \Add2~79\ ) + ( \Add2~78\ ))
-- \Add2~83\ = SHARE((!\R.aluData2\(20) & \R.aluData1\(20)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000010100000101000000000000000001010010110100101",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(20),
	datac => \ALT_INV_R.aluData1\(20),
	cin => \Add2~78\,
	sharein => \Add2~79\,
	sumout => \Add2~81_sumout\,
	cout => \Add2~82\,
	shareout => \Add2~83\);

-- Location: LABCELL_X79_Y5_N3
\Add2~85\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~85_sumout\ = SUM(( !\R.aluData1\(21) $ (\R.aluData2\(21)) ) + ( \Add2~83\ ) + ( \Add2~82\ ))
-- \Add2~86\ = CARRY(( !\R.aluData1\(21) $ (\R.aluData2\(21)) ) + ( \Add2~83\ ) + ( \Add2~82\ ))
-- \Add2~87\ = SHARE((\R.aluData1\(21) & !\R.aluData2\(21)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000000000000000000000001111000000001111",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluData1\(21),
	datad => \ALT_INV_R.aluData2\(21),
	cin => \Add2~82\,
	sharein => \Add2~83\,
	sumout => \Add2~85_sumout\,
	cout => \Add2~86\,
	shareout => \Add2~87\);

-- Location: LABCELL_X83_Y4_N15
\Selector13~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector13~3_combout\ = ( \Selector13~1_combout\ & ( (!\Selector13~0_combout\ & !\R.aluData2\(4)) ) ) # ( !\Selector13~1_combout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111111111111111111110100000101000001010000010100000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector13~0_combout\,
	datac => \ALT_INV_R.aluData2\(4),
	dataf => \ALT_INV_Selector13~1_combout\,
	combout => \Selector13~3_combout\);

-- Location: FF_X83_Y4_N16
\R.aluRes[19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector13~3_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(19));

-- Location: LABCELL_X77_Y9_N36
\Selector11~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector11~0_combout\ = ( \R.aluData2\(3) & ( \R.aluOp.ALUOpSRL~q\ & ( (\ShiftRight0~0_OTERM17\ & !\R.aluData2\(2)) ) ) ) # ( !\R.aluData2\(3) & ( \R.aluOp.ALUOpSRL~q\ & ( (!\R.aluData2\(2) & ((\ShiftRight1~11_OTERM35\))) # (\R.aluData2\(2) & 
-- (\ShiftRight1~12_OTERM57\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000110011010101010000111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~12_OTERM57\,
	datab => \ALT_INV_ShiftRight1~11_OTERM35\,
	datac => \ALT_INV_ShiftRight0~0_OTERM17\,
	datad => \ALT_INV_R.aluData2\(2),
	datae => \ALT_INV_R.aluData2\(3),
	dataf => \ALT_INV_R.aluOp.ALUOpSRL~q\,
	combout => \Selector11~0_combout\);

-- Location: LABCELL_X75_Y7_N18
\ShiftLeft0~12\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~12_combout\ = ( \Mux245~0_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (\Mux247~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & ((\Mux248~0_combout\))) ) ) ) # ( !\Mux245~0_combout\ & ( 
-- \NxR.aluData2[1]~17_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (\Mux247~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & ((\Mux248~0_combout\))) ) ) ) # ( \Mux245~0_combout\ & ( !\NxR.aluData2[1]~17_combout\ & ( (!\NxR.aluData2[0]~16_combout\) # 
-- (\Mux246~0_combout\) ) ) ) # ( !\Mux245~0_combout\ & ( !\NxR.aluData2[1]~17_combout\ & ( (\Mux246~0_combout\ & \NxR.aluData2[0]~16_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010101111111110101010100110011000011110011001100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux246~0_combout\,
	datab => \ALT_INV_Mux247~0_combout\,
	datac => \ALT_INV_Mux248~0_combout\,
	datad => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datae => \ALT_INV_Mux245~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[1]~17_combout\,
	combout => \ShiftLeft0~12_combout\);

-- Location: FF_X75_Y7_N19
\ShiftLeft0~12_NEW_REG790\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~12_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~12_OTERM791\);

-- Location: LABCELL_X73_Y6_N42
\ShiftLeft0~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~26_combout\ = ( \Mux238~0_combout\ & ( \NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\) # (\Mux240~0_combout\) ) ) ) # ( !\Mux238~0_combout\ & ( \NxR.aluData2[0]~16_combout\ & ( (\Mux240~0_combout\ & 
-- \NxR.aluData2[1]~17_combout\) ) ) ) # ( \Mux238~0_combout\ & ( !\NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (\Mux237~0_combout\)) # (\NxR.aluData2[1]~17_combout\ & ((\Mux239~0_combout\))) ) ) ) # ( !\Mux238~0_combout\ & ( 
-- !\NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (\Mux237~0_combout\)) # (\NxR.aluData2[1]~17_combout\ & ((\Mux239~0_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010100001111010101010000111100000000001100111111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux237~0_combout\,
	datab => \ALT_INV_Mux240~0_combout\,
	datac => \ALT_INV_Mux239~0_combout\,
	datad => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datae => \ALT_INV_Mux238~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[0]~16_combout\,
	combout => \ShiftLeft0~26_combout\);

-- Location: FF_X73_Y6_N43
\ShiftLeft0~26_NEW_REG738\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~26_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~26_OTERM739\);

-- Location: LABCELL_X74_Y6_N36
\ShiftLeft0~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~18_combout\ = ( \Mux243~0_combout\ & ( \Mux244~0_combout\ & ( ((!\NxR.aluData2[0]~16_combout\ & (\Mux241~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & ((\Mux242~0_combout\)))) # (\NxR.aluData2[1]~17_combout\) ) ) ) # ( !\Mux243~0_combout\ & ( 
-- \Mux244~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((!\NxR.aluData2[0]~16_combout\ & (\Mux241~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & ((\Mux242~0_combout\))))) # (\NxR.aluData2[1]~17_combout\ & (((\NxR.aluData2[0]~16_combout\)))) ) ) ) # ( 
-- \Mux243~0_combout\ & ( !\Mux244~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((!\NxR.aluData2[0]~16_combout\ & (\Mux241~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & ((\Mux242~0_combout\))))) # (\NxR.aluData2[1]~17_combout\ & 
-- (((!\NxR.aluData2[0]~16_combout\)))) ) ) ) # ( !\Mux243~0_combout\ & ( !\Mux244~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((!\NxR.aluData2[0]~16_combout\ & (\Mux241~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & ((\Mux242~0_combout\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010001000001010011101110000101000100010010111110111011101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datab => \ALT_INV_Mux241~0_combout\,
	datac => \ALT_INV_Mux242~0_combout\,
	datad => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datae => \ALT_INV_Mux243~0_combout\,
	dataf => \ALT_INV_Mux244~0_combout\,
	combout => \ShiftLeft0~18_combout\);

-- Location: FF_X74_Y6_N37
\ShiftLeft0~18_NEW_REG288\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~18_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~18_OTERM289\);

-- Location: LABCELL_X74_Y5_N48
\ShiftLeft0~34\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~34_combout\ = ( \NxR.aluData2[1]~17_combout\ & ( \Mux236~0_combout\ & ( (\Mux235~0_combout\) # (\NxR.aluData2[0]~16_combout\) ) ) ) # ( !\NxR.aluData2[1]~17_combout\ & ( \Mux236~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & 
-- (\Mux233~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & ((\Mux234~0_combout\))) ) ) ) # ( \NxR.aluData2[1]~17_combout\ & ( !\Mux236~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & \Mux235~0_combout\) ) ) ) # ( !\NxR.aluData2[1]~17_combout\ & ( 
-- !\Mux236~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (\Mux233~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & ((\Mux234~0_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101001101010011000000001111000001010011010100110000111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux233~0_combout\,
	datab => \ALT_INV_Mux234~0_combout\,
	datac => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datad => \ALT_INV_Mux235~0_combout\,
	datae => \ALT_INV_NxR.aluData2[1]~17_combout\,
	dataf => \ALT_INV_Mux236~0_combout\,
	combout => \ShiftLeft0~34_combout\);

-- Location: FF_X74_Y5_N49
\ShiftLeft0~34_NEW_REG298\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~34_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~34_OTERM299\);

-- Location: LABCELL_X77_Y9_N30
\ShiftLeft0~35\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~35_combout\ = ( \ShiftLeft0~18_OTERM289\ & ( \ShiftLeft0~34_OTERM299\ & ( (!\R.aluData2\(2)) # ((!\R.aluData2\(3) & ((\ShiftLeft0~26_OTERM739\))) # (\R.aluData2\(3) & (\ShiftLeft0~12_OTERM791\))) ) ) ) # ( !\ShiftLeft0~18_OTERM289\ & ( 
-- \ShiftLeft0~34_OTERM299\ & ( (!\R.aluData2\(3) & ((!\R.aluData2\(2)) # ((\ShiftLeft0~26_OTERM739\)))) # (\R.aluData2\(3) & (\R.aluData2\(2) & (\ShiftLeft0~12_OTERM791\))) ) ) ) # ( \ShiftLeft0~18_OTERM289\ & ( !\ShiftLeft0~34_OTERM299\ & ( 
-- (!\R.aluData2\(3) & (\R.aluData2\(2) & ((\ShiftLeft0~26_OTERM739\)))) # (\R.aluData2\(3) & ((!\R.aluData2\(2)) # ((\ShiftLeft0~12_OTERM791\)))) ) ) ) # ( !\ShiftLeft0~18_OTERM289\ & ( !\ShiftLeft0~34_OTERM299\ & ( (\R.aluData2\(2) & ((!\R.aluData2\(3) & 
-- ((\ShiftLeft0~26_OTERM739\))) # (\R.aluData2\(3) & (\ShiftLeft0~12_OTERM791\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000100100011010001010110011110001001101010111100110111101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(3),
	datab => \ALT_INV_R.aluData2\(2),
	datac => \ALT_INV_ShiftLeft0~12_OTERM791\,
	datad => \ALT_INV_ShiftLeft0~26_OTERM739\,
	datae => \ALT_INV_ShiftLeft0~18_OTERM289\,
	dataf => \ALT_INV_ShiftLeft0~34_OTERM299\,
	combout => \ShiftLeft0~35_combout\);

-- Location: LABCELL_X77_Y9_N24
\Selector11~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector11~1_combout\ = ( \R.aluOp.ALUOpSLL~q\ & ( \ShiftRight1~41_combout\ & ( (!\R.aluData2\(4) & (((\ShiftLeft0~35_combout\) # (\Selector11~0_combout\)) # (\R.aluOp.ALUOpSRA~q\))) ) ) ) # ( !\R.aluOp.ALUOpSLL~q\ & ( \ShiftRight1~41_combout\ & ( 
-- (!\R.aluData2\(4) & ((\Selector11~0_combout\) # (\R.aluOp.ALUOpSRA~q\))) ) ) ) # ( \R.aluOp.ALUOpSLL~q\ & ( !\ShiftRight1~41_combout\ & ( (!\R.aluData2\(4) & ((\ShiftLeft0~35_combout\) # (\Selector11~0_combout\))) ) ) ) # ( !\R.aluOp.ALUOpSLL~q\ & ( 
-- !\ShiftRight1~41_combout\ & ( (!\R.aluData2\(4) & \Selector11~0_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101000001010000010101010101000101010001010100010101010101010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(4),
	datab => \ALT_INV_R.aluOp.ALUOpSRA~q\,
	datac => \ALT_INV_Selector11~0_combout\,
	datad => \ALT_INV_ShiftLeft0~35_combout\,
	datae => \ALT_INV_R.aluOp.ALUOpSLL~q\,
	dataf => \ALT_INV_ShiftRight1~41_combout\,
	combout => \Selector11~1_combout\);

-- Location: FF_X78_Y2_N56
\R.aluRes[21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector11~5_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(21));

-- Location: MLABCELL_X78_Y5_N0
\Add1~81\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~81_sumout\ = SUM(( \R.aluData1\(20) ) + ( \R.aluData2\(20) ) + ( \Add1~78\ ))
-- \Add1~82\ = CARRY(( \R.aluData1\(20) ) + ( \R.aluData2\(20) ) + ( \Add1~78\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluData1\(20),
	dataf => \ALT_INV_R.aluData2\(20),
	cin => \Add1~78\,
	sumout => \Add1~81_sumout\,
	cout => \Add1~82\);

-- Location: MLABCELL_X78_Y5_N3
\Add1~85\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~85_sumout\ = SUM(( \R.aluData2\(21) ) + ( \R.aluData1\(21) ) + ( \Add1~82\ ))
-- \Add1~86\ = CARRY(( \R.aluData2\(21) ) + ( \R.aluData1\(21) ) + ( \Add1~82\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(21),
	datac => \ALT_INV_R.aluData1\(21),
	cin => \Add1~82\,
	sumout => \Add1~85_sumout\,
	cout => \Add1~86\);

-- Location: MLABCELL_X82_Y4_N42
\Equal3~5_RESYN1100\ : cyclonev_lcell_comb
-- Equation(s):
-- \Equal3~5_RESYN1100_BDD1101\ = ( \R.aluCalc~q\ & ( \Add1~85_sumout\ & ( (!\Selector11~1_combout\ & !\R.aluOp.ALUOpAdd~q\) ) ) ) # ( !\R.aluCalc~q\ & ( \Add1~85_sumout\ & ( (!\R.aluRes\(19) & !\R.aluRes\(21)) ) ) ) # ( \R.aluCalc~q\ & ( !\Add1~85_sumout\ & 
-- ( !\Selector11~1_combout\ ) ) ) # ( !\R.aluCalc~q\ & ( !\Add1~85_sumout\ & ( (!\R.aluRes\(19) & !\R.aluRes\(21)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010000010100000110011001100110010100000101000001100110000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluRes\(19),
	datab => \ALT_INV_Selector11~1_combout\,
	datac => \ALT_INV_R.aluRes\(21),
	datad => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datae => \ALT_INV_R.aluCalc~q\,
	dataf => \ALT_INV_Add1~85_sumout\,
	combout => \Equal3~5_RESYN1100_BDD1101\);

-- Location: LABCELL_X83_Y4_N12
\Equal3~5_RESYN1102\ : cyclonev_lcell_comb
-- Equation(s):
-- \Equal3~5_RESYN1102_BDD1103\ = (\Selector11~4_combout\ & !\Selector13~2_combout\)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100000000000011110000000000001111000000000000111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Selector11~4_combout\,
	datad => \ALT_INV_Selector13~2_combout\,
	combout => \Equal3~5_RESYN1102_BDD1103\);

-- Location: LABCELL_X83_Y4_N30
\Equal3~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Equal3~5_combout\ = ( \Equal3~5_RESYN1100_BDD1101\ & ( \Equal3~5_RESYN1102_BDD1103\ & ( (!\R.aluCalc~q\) # ((\Selector13~1_combout\ & ((!\R.aluOp.ALUOpSub~q\) # (!\Add2~85_sumout\)))) ) ) ) # ( \Equal3~5_RESYN1100_BDD1101\ & ( 
-- !\Equal3~5_RESYN1102_BDD1103\ & ( !\R.aluCalc~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000001111010111110100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector13~1_combout\,
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_R.aluCalc~q\,
	datad => \ALT_INV_Add2~85_sumout\,
	datae => \ALT_INV_Equal3~5_RESYN1100_BDD1101\,
	dataf => \ALT_INV_Equal3~5_RESYN1102_BDD1103\,
	combout => \Equal3~5_combout\);

-- Location: FF_X83_Y4_N31
\R.statusReg[0]_OTERM9_NEW_REG472\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Equal3~5_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.statusReg[0]_OTERM9_OTERM473\);

-- Location: LABCELL_X79_Y5_N6
\Add2~89\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~89_sumout\ = SUM(( !\R.aluData1\(22) $ (\R.aluData2\(22)) ) + ( \Add2~87\ ) + ( \Add2~86\ ))
-- \Add2~90\ = CARRY(( !\R.aluData1\(22) $ (\R.aluData2\(22)) ) + ( \Add2~87\ ) + ( \Add2~86\ ))
-- \Add2~91\ = SHARE((\R.aluData1\(22) & !\R.aluData2\(22)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000001100110000000000000000000000001100110000110011",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluData1\(22),
	datad => \ALT_INV_R.aluData2\(22),
	cin => \Add2~86\,
	sharein => \Add2~87\,
	sumout => \Add2~89_sumout\,
	cout => \Add2~90\,
	shareout => \Add2~91\);

-- Location: LABCELL_X79_Y5_N9
\Add2~93\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~93_sumout\ = SUM(( !\R.aluData1\(23) $ (\R.aluData2\(23)) ) + ( \Add2~91\ ) + ( \Add2~90\ ))
-- \Add2~94\ = CARRY(( !\R.aluData1\(23) $ (\R.aluData2\(23)) ) + ( \Add2~91\ ) + ( \Add2~90\ ))
-- \Add2~95\ = SHARE((\R.aluData1\(23) & !\R.aluData2\(23)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010101010000000000000000000000001010101001010101",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData1\(23),
	datad => \ALT_INV_R.aluData2\(23),
	cin => \Add2~90\,
	sharein => \Add2~91\,
	sumout => \Add2~93_sumout\,
	cout => \Add2~94\,
	shareout => \Add2~95\);

-- Location: LABCELL_X79_Y5_N12
\Add2~97\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~97_sumout\ = SUM(( !\R.aluData2\(24) $ (\R.aluData1\(24)) ) + ( \Add2~95\ ) + ( \Add2~94\ ))
-- \Add2~98\ = CARRY(( !\R.aluData2\(24) $ (\R.aluData1\(24)) ) + ( \Add2~95\ ) + ( \Add2~94\ ))
-- \Add2~99\ = SHARE((!\R.aluData2\(24) & \R.aluData1\(24)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011000000110000000000000000001100001111000011",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluData2\(24),
	datac => \ALT_INV_R.aluData1\(24),
	cin => \Add2~94\,
	sharein => \Add2~95\,
	sumout => \Add2~97_sumout\,
	cout => \Add2~98\,
	shareout => \Add2~99\);

-- Location: LABCELL_X79_Y5_N15
\Add2~101\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~101_sumout\ = SUM(( !\R.aluData1\(25) $ (\R.aluData2[25]~DUPLICATE_q\) ) + ( \Add2~99\ ) + ( \Add2~98\ ))
-- \Add2~102\ = CARRY(( !\R.aluData1\(25) $ (\R.aluData2[25]~DUPLICATE_q\) ) + ( \Add2~99\ ) + ( \Add2~98\ ))
-- \Add2~103\ = SHARE((\R.aluData1\(25) & !\R.aluData2[25]~DUPLICATE_q\))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010101010000000000000000000000001010101001010101",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData1\(25),
	datad => \ALT_INV_R.aluData2[25]~DUPLICATE_q\,
	cin => \Add2~98\,
	sharein => \Add2~99\,
	sumout => \Add2~101_sumout\,
	cout => \Add2~102\,
	shareout => \Add2~103\);

-- Location: LABCELL_X79_Y5_N18
\Add2~105\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~105_sumout\ = SUM(( !\R.aluData2\(26) $ (\R.aluData1\(26)) ) + ( \Add2~103\ ) + ( \Add2~102\ ))
-- \Add2~106\ = CARRY(( !\R.aluData2\(26) $ (\R.aluData1\(26)) ) + ( \Add2~103\ ) + ( \Add2~102\ ))
-- \Add2~107\ = SHARE((!\R.aluData2\(26) & \R.aluData1\(26)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011000000110000000000000000001100001111000011",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluData2\(26),
	datac => \ALT_INV_R.aluData1\(26),
	cin => \Add2~102\,
	sharein => \Add2~103\,
	sumout => \Add2~105_sumout\,
	cout => \Add2~106\,
	shareout => \Add2~107\);

-- Location: LABCELL_X79_Y5_N21
\Add2~109\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~109_sumout\ = SUM(( !\R.aluData1\(27) $ (\R.aluData2\(27)) ) + ( \Add2~107\ ) + ( \Add2~106\ ))
-- \Add2~110\ = CARRY(( !\R.aluData1\(27) $ (\R.aluData2\(27)) ) + ( \Add2~107\ ) + ( \Add2~106\ ))
-- \Add2~111\ = SHARE((\R.aluData1\(27) & !\R.aluData2\(27)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010100000101000000000000000000001010010110100101",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData1\(27),
	datac => \ALT_INV_R.aluData2\(27),
	cin => \Add2~106\,
	sharein => \Add2~107\,
	sumout => \Add2~109_sumout\,
	cout => \Add2~110\,
	shareout => \Add2~111\);

-- Location: LABCELL_X74_Y3_N54
\ShiftLeft0~38\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~38_combout\ = ( \NxR.aluData2[0]~16_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( \Mux234~0_combout\ ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( \Mux233~0_combout\ ) ) ) # ( \NxR.aluData2[0]~16_combout\ & ( 
-- !\NxR.aluData2[1]~17_combout\ & ( \Mux232~0_combout\ ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( !\NxR.aluData2[1]~17_combout\ & ( \Mux231~0_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110011010101010101010100001111000011110000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux232~0_combout\,
	datab => \ALT_INV_Mux231~0_combout\,
	datac => \ALT_INV_Mux233~0_combout\,
	datad => \ALT_INV_Mux234~0_combout\,
	datae => \ALT_INV_NxR.aluData2[0]~16_combout\,
	dataf => \ALT_INV_NxR.aluData2[1]~17_combout\,
	combout => \ShiftLeft0~38_combout\);

-- Location: FF_X74_Y3_N55
\ShiftLeft0~38_NEW_REG788\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~38_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~38_OTERM789\);

-- Location: LABCELL_X73_Y4_N30
\ShiftLeft0~47\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~47_combout\ = ( \Mux227~0_combout\ & ( \Mux229~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\) # ((!\NxR.aluData2[1]~17_combout\ & (\Mux228~0_combout\)) # (\NxR.aluData2[1]~17_combout\ & ((\Mux230~0_combout\)))) ) ) ) # ( !\Mux227~0_combout\ & 
-- ( \Mux229~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (((\NxR.aluData2[1]~17_combout\)))) # (\NxR.aluData2[0]~16_combout\ & ((!\NxR.aluData2[1]~17_combout\ & (\Mux228~0_combout\)) # (\NxR.aluData2[1]~17_combout\ & ((\Mux230~0_combout\))))) ) ) ) # ( 
-- \Mux227~0_combout\ & ( !\Mux229~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (((!\NxR.aluData2[1]~17_combout\)))) # (\NxR.aluData2[0]~16_combout\ & ((!\NxR.aluData2[1]~17_combout\ & (\Mux228~0_combout\)) # (\NxR.aluData2[1]~17_combout\ & 
-- ((\Mux230~0_combout\))))) ) ) ) # ( !\Mux227~0_combout\ & ( !\Mux229~0_combout\ & ( (\NxR.aluData2[0]~16_combout\ & ((!\NxR.aluData2[1]~17_combout\ & (\Mux228~0_combout\)) # (\NxR.aluData2[1]~17_combout\ & ((\Mux230~0_combout\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000000010101101100001011010100011010000111111011101010111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datab => \ALT_INV_Mux228~0_combout\,
	datac => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datad => \ALT_INV_Mux230~0_combout\,
	datae => \ALT_INV_Mux227~0_combout\,
	dataf => \ALT_INV_Mux229~0_combout\,
	combout => \ShiftLeft0~47_combout\);

-- Location: FF_X73_Y4_N31
\ShiftLeft0~47_NEW_REG758\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~47_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~47_OTERM759\);

-- Location: LABCELL_X74_Y6_N18
\ShiftLeft0~30\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~30_combout\ = ( \Mux238~0_combout\ & ( \NxR.aluData2[0]~16_combout\ & ( (\Mux236~0_combout\) # (\NxR.aluData2[1]~17_combout\) ) ) ) # ( !\Mux238~0_combout\ & ( \NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & 
-- \Mux236~0_combout\) ) ) ) # ( \Mux238~0_combout\ & ( !\NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((\Mux235~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux237~0_combout\)) ) ) ) # ( !\Mux238~0_combout\ & ( 
-- !\NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((\Mux235~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux237~0_combout\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010110101111000001011010111100100010001000100111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datab => \ALT_INV_Mux236~0_combout\,
	datac => \ALT_INV_Mux237~0_combout\,
	datad => \ALT_INV_Mux235~0_combout\,
	datae => \ALT_INV_Mux238~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[0]~16_combout\,
	combout => \ShiftLeft0~30_combout\);

-- Location: FF_X74_Y6_N19
\ShiftLeft0~30_NEW_REG600\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~30_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~30_OTERM601\);

-- Location: LABCELL_X73_Y8_N48
\ShiftLeft0~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~22_combout\ = ( \Mux241~0_combout\ & ( \NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((\Mux240~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux242~0_combout\)) ) ) ) # ( !\Mux241~0_combout\ & ( 
-- \NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((\Mux240~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux242~0_combout\)) ) ) ) # ( \Mux241~0_combout\ & ( !\NxR.aluData2[0]~16_combout\ & ( (\Mux239~0_combout\) # 
-- (\NxR.aluData2[1]~17_combout\) ) ) ) # ( !\Mux241~0_combout\ & ( !\NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & \Mux239~0_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101000001010010111110101111100010001101110110001000110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datab => \ALT_INV_Mux242~0_combout\,
	datac => \ALT_INV_Mux239~0_combout\,
	datad => \ALT_INV_Mux240~0_combout\,
	datae => \ALT_INV_Mux241~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[0]~16_combout\,
	combout => \ShiftLeft0~22_combout\);

-- Location: FF_X73_Y8_N49
\ShiftLeft0~22_NEW_REG736\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~22_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~22_OTERM737\);

-- Location: LABCELL_X79_Y7_N48
\ShiftLeft0~48\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~48_combout\ = ( \ShiftLeft0~22_OTERM737\ & ( \R.aluData2\(2) & ( (\R.aluData2\(3)) # (\ShiftLeft0~38_OTERM789\) ) ) ) # ( !\ShiftLeft0~22_OTERM737\ & ( \R.aluData2\(2) & ( (\ShiftLeft0~38_OTERM789\ & !\R.aluData2\(3)) ) ) ) # ( 
-- \ShiftLeft0~22_OTERM737\ & ( !\R.aluData2\(2) & ( (!\R.aluData2\(3) & (\ShiftLeft0~47_OTERM759\)) # (\R.aluData2\(3) & ((\ShiftLeft0~30_OTERM601\))) ) ) ) # ( !\ShiftLeft0~22_OTERM737\ & ( !\R.aluData2\(2) & ( (!\R.aluData2\(3) & 
-- (\ShiftLeft0~47_OTERM759\)) # (\R.aluData2\(3) & ((\ShiftLeft0~30_OTERM601\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100001111001100110000111101010101000000000101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~38_OTERM789\,
	datab => \ALT_INV_ShiftLeft0~47_OTERM759\,
	datac => \ALT_INV_ShiftLeft0~30_OTERM601\,
	datad => \ALT_INV_R.aluData2\(3),
	datae => \ALT_INV_ShiftLeft0~22_OTERM737\,
	dataf => \ALT_INV_R.aluData2\(2),
	combout => \ShiftLeft0~48_combout\);

-- Location: LABCELL_X73_Y5_N12
\ShiftRight1~32\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~32_combout\ = ( \NxR.aluData2[0]~16_combout\ & ( \Mux226~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\) # (\Mux224~0_combout\) ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( \Mux226~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & 
-- ((\Mux227~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux225~0_combout\)) ) ) ) # ( \NxR.aluData2[0]~16_combout\ & ( !\Mux226~0_combout\ & ( (\Mux224~0_combout\ & \NxR.aluData2[1]~17_combout\) ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( 
-- !\Mux226~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((\Mux227~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux225~0_combout\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111101010101000000000011001100001111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux225~0_combout\,
	datab => \ALT_INV_Mux224~0_combout\,
	datac => \ALT_INV_Mux227~0_combout\,
	datad => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datae => \ALT_INV_NxR.aluData2[0]~16_combout\,
	dataf => \ALT_INV_Mux226~0_combout\,
	combout => \ShiftRight1~32_combout\);

-- Location: FF_X73_Y5_N13
\ShiftRight1~32_NEW_REG20\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~32_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~32_OTERM21\);

-- Location: LABCELL_X73_Y6_N39
\ShiftRight0~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight0~4_combout\ = ( !\NxR.aluData2[0]~16_combout\ & ( (\Mux223~0_combout\ & !\NxR.aluData2[1]~17_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100000000000011110000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Mux223~0_combout\,
	datad => \ALT_INV_NxR.aluData2[1]~17_combout\,
	dataf => \ALT_INV_NxR.aluData2[0]~16_combout\,
	combout => \ShiftRight0~4_combout\);

-- Location: FF_X73_Y6_N41
\ShiftRight0~4_NEW_REG30\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight0~4_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight0~4_OTERM31\);

-- Location: LABCELL_X79_Y7_N45
\Selector5~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector5~0_combout\ = ( \R.aluOp.ALUOpSRL~q\ & ( (!\R.aluData2\(3) & ((!\R.aluData2\(2) & (\ShiftRight1~32_OTERM21\)) # (\R.aluData2\(2) & ((\ShiftRight0~4_OTERM31\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000001000111000000000100011100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~32_OTERM21\,
	datab => \ALT_INV_R.aluData2\(2),
	datac => \ALT_INV_ShiftRight0~4_OTERM31\,
	datad => \ALT_INV_R.aluData2\(3),
	dataf => \ALT_INV_R.aluOp.ALUOpSRL~q\,
	combout => \Selector5~0_combout\);

-- Location: LABCELL_X79_Y7_N42
\Selector5~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector5~1_combout\ = ( \ShiftRight0~7_OTERM233DUPLICATE_q\ & ( (\R.aluData1\(31) & \R.aluOp.ALUOpSRA~q\) ) ) # ( !\ShiftRight0~7_OTERM233DUPLICATE_q\ & ( (\ShiftRight1~32_OTERM21\ & \R.aluOp.ALUOpSRA~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010101000000000101010100000000000011110000000000001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~32_OTERM21\,
	datac => \ALT_INV_R.aluData1\(31),
	datad => \ALT_INV_R.aluOp.ALUOpSRA~q\,
	dataf => \ALT_INV_ShiftRight0~7_OTERM233DUPLICATE_q\,
	combout => \Selector5~1_combout\);

-- Location: LABCELL_X79_Y7_N6
\Selector5~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector5~2_combout\ = ( \Selector5~0_combout\ & ( \Selector5~1_combout\ & ( !\R.aluData2\(4) ) ) ) # ( !\Selector5~0_combout\ & ( \Selector5~1_combout\ & ( !\R.aluData2\(4) ) ) ) # ( \Selector5~0_combout\ & ( !\Selector5~1_combout\ & ( !\R.aluData2\(4) 
-- ) ) ) # ( !\Selector5~0_combout\ & ( !\Selector5~1_combout\ & ( (\ShiftLeft0~48_combout\ & (!\R.aluData2\(4) & \R.aluOp.ALUOpSLL~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010000111100001111000011110000111100001111000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~48_combout\,
	datac => \ALT_INV_R.aluData2\(4),
	datad => \ALT_INV_R.aluOp.ALUOpSLL~q\,
	datae => \ALT_INV_Selector5~0_combout\,
	dataf => \ALT_INV_Selector5~1_combout\,
	combout => \Selector5~2_combout\);

-- Location: LABCELL_X74_Y7_N48
\ShiftLeft0~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~9_combout\ = ( \Mux247~0_combout\ & ( \Mux250~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((!\NxR.aluData2[0]~16_combout\) # (\Mux248~0_combout\)))) # (\NxR.aluData2[1]~17_combout\ & (((\NxR.aluData2[0]~16_combout\)) # 
-- (\Mux249~0_combout\))) ) ) ) # ( !\Mux247~0_combout\ & ( \Mux250~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((\Mux248~0_combout\ & \NxR.aluData2[0]~16_combout\)))) # (\NxR.aluData2[1]~17_combout\ & (((\NxR.aluData2[0]~16_combout\)) # 
-- (\Mux249~0_combout\))) ) ) ) # ( \Mux247~0_combout\ & ( !\Mux250~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((!\NxR.aluData2[0]~16_combout\) # (\Mux248~0_combout\)))) # (\NxR.aluData2[1]~17_combout\ & (\Mux249~0_combout\ & 
-- ((!\NxR.aluData2[0]~16_combout\)))) ) ) ) # ( !\Mux247~0_combout\ & ( !\Mux250~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((\Mux248~0_combout\ & \NxR.aluData2[0]~16_combout\)))) # (\NxR.aluData2[1]~17_combout\ & (\Mux249~0_combout\ & 
-- ((!\NxR.aluData2[0]~16_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100001100110111010000110000010001001111111101110100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux249~0_combout\,
	datab => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datac => \ALT_INV_Mux248~0_combout\,
	datad => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datae => \ALT_INV_Mux247~0_combout\,
	dataf => \ALT_INV_Mux250~0_combout\,
	combout => \ShiftLeft0~9_combout\);

-- Location: FF_X74_Y7_N49
\ShiftLeft0~9_NEW_REG460\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~9_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~9_OTERM461\);

-- Location: LABCELL_X77_Y8_N21
\ShiftLeft0~15\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~15_combout\ = ( \ShiftLeft0~9_OTERM461\ & ( (!\R.aluData2\(3) & (((\ShiftLeft0~14_OTERM753\)) # (\R.aluData2\(2)))) # (\R.aluData2\(3) & (!\R.aluData2\(2) & (\ShiftLeft0~3_OTERM223\))) ) ) # ( !\ShiftLeft0~9_OTERM461\ & ( (!\R.aluData2\(2) & 
-- ((!\R.aluData2\(3) & ((\ShiftLeft0~14_OTERM753\))) # (\R.aluData2\(3) & (\ShiftLeft0~3_OTERM223\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010010001100000001001000110000100110101011100010011010101110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(3),
	datab => \ALT_INV_R.aluData2\(2),
	datac => \ALT_INV_ShiftLeft0~3_OTERM223\,
	datad => \ALT_INV_ShiftLeft0~14_OTERM753\,
	dataf => \ALT_INV_ShiftLeft0~9_OTERM461\,
	combout => \ShiftLeft0~15_combout\);

-- Location: LABCELL_X77_Y8_N6
\Selector5~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector5~3_combout\ = ( \R.aluData1\(27) & ( (!\R.aluOp.ALUOpOr~q\ & ((!\R.aluData2\(27) & ((!\R.aluOp.ALUOpXor~DUPLICATE_q\))) # (\R.aluData2\(27) & (!\R.aluOp.ALUOpAnd~DUPLICATE_q\)))) ) ) # ( !\R.aluData1\(27) & ( (!\R.aluData2\(27)) # 
-- ((!\R.aluOp.ALUOpOr~q\ & !\R.aluOp.ALUOpXor~DUPLICATE_q\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111110011110000111111001111000011001000000010001100100000001000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpAnd~DUPLICATE_q\,
	datab => \ALT_INV_R.aluOp.ALUOpOr~q\,
	datac => \ALT_INV_R.aluData2\(27),
	datad => \ALT_INV_R.aluOp.ALUOpXor~DUPLICATE_q\,
	dataf => \ALT_INV_R.aluData1\(27),
	combout => \Selector5~3_combout\);

-- Location: LABCELL_X77_Y8_N3
\Selector5~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector5~4_combout\ = ( \Selector5~3_combout\ & ( (!\Selector17~0_OTERM391\ & ((!\ShiftLeft0~15_combout\) # (!\Selector12~2_OTERM395\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000010101010101000001010101010100000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector17~0_OTERM391\,
	datac => \ALT_INV_ShiftLeft0~15_combout\,
	datad => \ALT_INV_Selector12~2_OTERM395\,
	dataf => \ALT_INV_Selector5~3_combout\,
	combout => \Selector5~4_combout\);

-- Location: LABCELL_X79_Y4_N12
\Selector5~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector5~5_combout\ = ( \Add1~109_sumout\ & ( \Add2~109_sumout\ & ( (((!\Selector5~4_combout\) # (\Selector5~2_combout\)) # (\R.aluOp.ALUOpSub~q\)) # (\R.aluOp.ALUOpAdd~q\) ) ) ) # ( !\Add1~109_sumout\ & ( \Add2~109_sumout\ & ( ((!\Selector5~4_combout\) 
-- # (\Selector5~2_combout\)) # (\R.aluOp.ALUOpSub~q\) ) ) ) # ( \Add1~109_sumout\ & ( !\Add2~109_sumout\ & ( ((!\Selector5~4_combout\) # (\Selector5~2_combout\)) # (\R.aluOp.ALUOpAdd~q\) ) ) ) # ( !\Add1~109_sumout\ & ( !\Add2~109_sumout\ & ( 
-- (!\Selector5~4_combout\) # (\Selector5~2_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111000011111111111101011111111111110011111111111111011111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_Selector5~4_combout\,
	datad => \ALT_INV_Selector5~2_combout\,
	datae => \ALT_INV_Add1~109_sumout\,
	dataf => \ALT_INV_Add2~109_sumout\,
	combout => \Selector5~5_combout\);

-- Location: FF_X79_Y4_N14
\R.aluRes[27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector5~5_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(27));

-- Location: LABCELL_X79_Y4_N45
\vAluRes~35\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~35_combout\ = ( \R.aluCalc~q\ & ( (!\Selector5~2_combout\ & \Selector5~4_combout\) ) ) # ( !\R.aluCalc~q\ & ( !\R.aluRes\(27) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111000011110000111100001111000000000000110011000000000011001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Selector5~2_combout\,
	datac => \ALT_INV_R.aluRes\(27),
	datad => \ALT_INV_Selector5~4_combout\,
	dataf => \ALT_INV_R.aluCalc~q\,
	combout => \vAluRes~35_combout\);

-- Location: LABCELL_X79_Y4_N6
\vAluRes~24\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~24_combout\ = ( \vAluRes~35_combout\ & ( \R.aluCalc~q\ & ( (!\R.aluOp.ALUOpAdd~q\ & (\Add2~109_sumout\ & ((\R.aluOp.ALUOpSub~q\)))) # (\R.aluOp.ALUOpAdd~q\ & (((\Add2~109_sumout\ & \R.aluOp.ALUOpSub~q\)) # (\Add1~109_sumout\))) ) ) ) # ( 
-- !\vAluRes~35_combout\ & ( \R.aluCalc~q\ ) ) # ( !\vAluRes~35_combout\ & ( !\R.aluCalc~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111000000000000000011111111111111110000010100110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datab => \ALT_INV_Add2~109_sumout\,
	datac => \ALT_INV_Add1~109_sumout\,
	datad => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datae => \ALT_INV_vAluRes~35_combout\,
	dataf => \ALT_INV_R.aluCalc~q\,
	combout => \vAluRes~24_combout\);

-- Location: FF_X79_Y4_N8
\R.statusReg[0]_OTERM9_NEW_REG466\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \vAluRes~24_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.statusReg[0]_OTERM9_OTERM467\);

-- Location: FF_X78_Y3_N56
\R.aluRes[17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector15~5_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(17));

-- Location: MLABCELL_X78_Y3_N12
\Equal3~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Equal3~14_combout\ = ( \Add1~65_sumout\ & ( \R.aluOp.ALUOpAdd~q\ & ( (!\R.aluRes\(16) & (!\R.aluRes\(17) & !\R.aluCalc~q\)) ) ) ) # ( !\Add1~65_sumout\ & ( \R.aluOp.ALUOpAdd~q\ & ( (!\R.aluCalc~q\ & (!\R.aluRes\(16) & ((!\R.aluRes\(17))))) # 
-- (\R.aluCalc~q\ & (((!\Add1~69_sumout\)))) ) ) ) # ( \Add1~65_sumout\ & ( !\R.aluOp.ALUOpAdd~q\ & ( ((!\R.aluRes\(16) & !\R.aluRes\(17))) # (\R.aluCalc~q\) ) ) ) # ( !\Add1~65_sumout\ & ( !\R.aluOp.ALUOpAdd~q\ & ( ((!\R.aluRes\(16) & !\R.aluRes\(17))) # 
-- (\R.aluCalc~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010000011111111101000001111111110100000110011001010000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluRes\(16),
	datab => \ALT_INV_Add1~69_sumout\,
	datac => \ALT_INV_R.aluRes\(17),
	datad => \ALT_INV_R.aluCalc~q\,
	datae => \ALT_INV_Add1~65_sumout\,
	dataf => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	combout => \Equal3~14_combout\);

-- Location: MLABCELL_X72_Y7_N3
\ShiftLeft0~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~1_combout\ = ( \NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & \Mux254~0_combout\) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( (\Mux253~0_combout\ & !\NxR.aluData2[1]~17_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101000001010000010100000101000000000000111100000000000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux253~0_combout\,
	datac => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datad => \ALT_INV_Mux254~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[0]~16_combout\,
	combout => \ShiftLeft0~1_combout\);

-- Location: FF_X72_Y7_N4
\ShiftLeft0~1_NEW_REG254\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~1_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~1_OTERM255\);

-- Location: MLABCELL_X72_Y5_N9
\Selector15~2_RTM0743\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector15~2_RTM0743_combout\ = ( \Mux237~0_combout\ & ( ((!\NxR.aluData2[17]~4_combout\ & (\R.aluOp.ALUOpXor_OTERM355\)) # (\NxR.aluData2[17]~4_combout\ & ((\R.aluOp.ALUOpAnd_OTERM357\)))) # (\R.aluOp.ALUOpOr_OTERM353\) ) ) # ( !\Mux237~0_combout\ & ( 
-- (\NxR.aluData2[17]~4_combout\ & ((\R.aluOp.ALUOpXor_OTERM355\) # (\R.aluOp.ALUOpOr_OTERM353\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001110111000000000111011101110111010111110111011101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpOr_OTERM353\,
	datab => \ALT_INV_R.aluOp.ALUOpXor_OTERM355\,
	datac => \ALT_INV_R.aluOp.ALUOpAnd_OTERM357\,
	datad => \ALT_INV_NxR.aluData2[17]~4_combout\,
	dataf => \ALT_INV_Mux237~0_combout\,
	combout => \Selector15~2_RTM0743_combout\);

-- Location: FF_X72_Y5_N10
\Selector15~2_NEW_REG740\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector15~2_RTM0743_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector15~2_OTERM741\);

-- Location: LABCELL_X73_Y7_N39
\Selector15~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector15~3_combout\ = (!\Selector15~2_OTERM741\ & ((!\Selector16~0_OTERM393\) # (!\ShiftLeft0~1_OTERM255\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111101000000000111110100000000011111010000000001111101000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector16~0_OTERM393\,
	datac => \ALT_INV_ShiftLeft0~1_OTERM255\,
	datad => \ALT_INV_Selector15~2_OTERM741\,
	combout => \Selector15~3_combout\);

-- Location: MLABCELL_X84_Y7_N24
\ShiftLeft0~27\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~27_combout\ = ( \ShiftLeft0~26_OTERM739\ & ( \R.aluData2\(2) & ( (!\R.aluData2\(3) & ((\ShiftLeft0~18_OTERM289\))) # (\R.aluData2\(3) & (\ShiftLeft0~7_OTERM205\)) ) ) ) # ( !\ShiftLeft0~26_OTERM739\ & ( \R.aluData2\(2) & ( (!\R.aluData2\(3) & 
-- ((\ShiftLeft0~18_OTERM289\))) # (\R.aluData2\(3) & (\ShiftLeft0~7_OTERM205\)) ) ) ) # ( \ShiftLeft0~26_OTERM739\ & ( !\R.aluData2\(2) & ( (!\R.aluData2\(3)) # (\ShiftLeft0~12_OTERM791\) ) ) ) # ( !\ShiftLeft0~26_OTERM739\ & ( !\R.aluData2\(2) & ( 
-- (\R.aluData2\(3) & \ShiftLeft0~12_OTERM791\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011110011111100111100010001110111010001000111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~7_OTERM205\,
	datab => \ALT_INV_R.aluData2\(3),
	datac => \ALT_INV_ShiftLeft0~12_OTERM791\,
	datad => \ALT_INV_ShiftLeft0~18_OTERM289\,
	datae => \ALT_INV_ShiftLeft0~26_OTERM739\,
	dataf => \ALT_INV_R.aluData2\(2),
	combout => \ShiftLeft0~27_combout\);

-- Location: LABCELL_X80_Y3_N6
\Selector15~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector15~4_combout\ = ( \R.aluOp.ALUOpSLL~q\ & ( \ShiftLeft0~27_combout\ & ( (\Selector15~3_combout\ & \R.aluData2\(4)) ) ) ) # ( !\R.aluOp.ALUOpSLL~q\ & ( \ShiftLeft0~27_combout\ & ( (\Selector15~3_combout\ & ((!\R.aluOp.ALUOpSRL~q\) # 
-- ((!\ShiftRight0~1_combout\) # (\R.aluData2\(4))))) ) ) ) # ( \R.aluOp.ALUOpSLL~q\ & ( !\ShiftLeft0~27_combout\ & ( (\Selector15~3_combout\ & ((!\R.aluOp.ALUOpSRL~q\) # ((!\ShiftRight0~1_combout\) # (\R.aluData2\(4))))) ) ) ) # ( !\R.aluOp.ALUOpSLL~q\ & ( 
-- !\ShiftLeft0~27_combout\ & ( (\Selector15~3_combout\ & ((!\R.aluOp.ALUOpSRL~q\) # ((!\ShiftRight0~1_combout\) # (\R.aluData2\(4))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010001010101010101000101010101010100010101010000000001010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector15~3_combout\,
	datab => \ALT_INV_R.aluOp.ALUOpSRL~q\,
	datac => \ALT_INV_ShiftRight0~1_combout\,
	datad => \ALT_INV_R.aluData2\(4),
	datae => \ALT_INV_R.aluOp.ALUOpSLL~q\,
	dataf => \ALT_INV_ShiftLeft0~27_combout\,
	combout => \Selector15~4_combout\);

-- Location: LABCELL_X77_Y9_N0
\ShiftRight1~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~14_combout\ = ( \R.aluData2\(3) & ( \ShiftRight1~13_OTERM15\ & ( (\R.aluData2\(2)) # (\ShiftRight1~12_OTERM57\) ) ) ) # ( !\R.aluData2\(3) & ( \ShiftRight1~13_OTERM15\ & ( (!\R.aluData2\(2) & (\ShiftRight1~10_OTERM265\)) # (\R.aluData2\(2) & 
-- ((\ShiftRight1~11_OTERM35\))) ) ) ) # ( \R.aluData2\(3) & ( !\ShiftRight1~13_OTERM15\ & ( (\ShiftRight1~12_OTERM57\ & !\R.aluData2\(2)) ) ) ) # ( !\R.aluData2\(3) & ( !\ShiftRight1~13_OTERM15\ & ( (!\R.aluData2\(2) & (\ShiftRight1~10_OTERM265\)) # 
-- (\R.aluData2\(2) & ((\ShiftRight1~11_OTERM35\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000110000111111010001000100010000001100001111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~12_OTERM57\,
	datab => \ALT_INV_R.aluData2\(2),
	datac => \ALT_INV_ShiftRight1~10_OTERM265\,
	datad => \ALT_INV_ShiftRight1~11_OTERM35\,
	datae => \ALT_INV_R.aluData2\(3),
	dataf => \ALT_INV_ShiftRight1~13_OTERM15\,
	combout => \ShiftRight1~14_combout\);

-- Location: LABCELL_X77_Y9_N45
\Selector15~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector15~0_combout\ = ( \R.aluData1\(31) & ( (\R.aluOp.ALUOpSRA~q\ & ((\ShiftRight1~14_combout\) # (\R.aluData2\(4)))) ) ) # ( !\R.aluData1\(31) & ( (!\R.aluData2\(4) & (\R.aluOp.ALUOpSRA~q\ & \ShiftRight1~14_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000001010000000000000101000000101000011110000010100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(4),
	datac => \ALT_INV_R.aluOp.ALUOpSRA~q\,
	datad => \ALT_INV_ShiftRight1~14_combout\,
	dataf => \ALT_INV_R.aluData1\(31),
	combout => \Selector15~0_combout\);

-- Location: MLABCELL_X78_Y3_N0
\Equal3~15\ : cyclonev_lcell_comb
-- Equation(s):
-- \Equal3~15_combout\ = (\Selector16~3_combout\ & (\Selector15~4_combout\ & !\Selector15~0_combout\))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100000000000100010000000000010001000000000001000100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector16~3_combout\,
	datab => \ALT_INV_Selector15~4_combout\,
	datad => \ALT_INV_Selector15~0_combout\,
	combout => \Equal3~15_combout\);

-- Location: LABCELL_X79_Y3_N18
\Equal3~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Equal3~4_combout\ = ( \R.aluOp.ALUOpSub~q\ & ( \Equal3~15_combout\ & ( (\Equal3~14_combout\ & ((!\R.aluCalc~q\) # ((!\Add2~69_sumout\ & !\Add2~65_sumout\)))) ) ) ) # ( !\R.aluOp.ALUOpSub~q\ & ( \Equal3~15_combout\ & ( \Equal3~14_combout\ ) ) ) # ( 
-- \R.aluOp.ALUOpSub~q\ & ( !\Equal3~15_combout\ & ( (\Equal3~14_combout\ & !\R.aluCalc~q\) ) ) ) # ( !\R.aluOp.ALUOpSub~q\ & ( !\Equal3~15_combout\ & ( (\Equal3~14_combout\ & !\R.aluCalc~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100010001000100010001000100010001010101010101010101010001000100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Equal3~14_combout\,
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_Add2~69_sumout\,
	datad => \ALT_INV_Add2~65_sumout\,
	datae => \ALT_INV_R.aluOp.ALUOpSub~q\,
	dataf => \ALT_INV_Equal3~15_combout\,
	combout => \Equal3~4_combout\);

-- Location: FF_X79_Y3_N19
\R.statusReg[0]_OTERM9_NEW_REG470\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Equal3~4_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.statusReg[0]_OTERM9_OTERM471\);

-- Location: FF_X83_Y6_N13
\R.statusReg[0]_OTERM9_NEW_REG462\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \vAluRes~60_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.statusReg[0]_OTERM9_OTERM463\);

-- Location: LABCELL_X73_Y8_N39
\ShiftLeft0~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~0_combout\ = ( !\NxR.aluData2[1]~17_combout\ & ( !\NxR.aluData2[0]~16_combout\ & ( \Mux254~0_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \ALT_INV_Mux254~0_combout\,
	datae => \ALT_INV_NxR.aluData2[1]~17_combout\,
	dataf => \ALT_INV_NxR.aluData2[0]~16_combout\,
	combout => \ShiftLeft0~0_combout\);

-- Location: FF_X73_Y8_N40
\ShiftLeft0~0_NEW_REG262\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~0_OTERM263\);

-- Location: LABCELL_X75_Y7_N48
\ShiftLeft0~16\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~16_combout\ = ( \Mux244~0_combout\ & ( \Mux243~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((\NxR.aluData2[0]~16_combout\)) # (\Mux242~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (((!\NxR.aluData2[0]~16_combout\) # 
-- (\Mux245~0_combout\)))) ) ) ) # ( !\Mux244~0_combout\ & ( \Mux243~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((\NxR.aluData2[0]~16_combout\)) # (\Mux242~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (((\NxR.aluData2[0]~16_combout\ & 
-- \Mux245~0_combout\)))) ) ) ) # ( \Mux244~0_combout\ & ( !\Mux243~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (\Mux242~0_combout\ & (!\NxR.aluData2[0]~16_combout\))) # (\NxR.aluData2[1]~17_combout\ & (((!\NxR.aluData2[0]~16_combout\) # 
-- (\Mux245~0_combout\)))) ) ) ) # ( !\Mux244~0_combout\ & ( !\Mux243~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (\Mux242~0_combout\ & (!\NxR.aluData2[0]~16_combout\))) # (\NxR.aluData2[1]~17_combout\ & (((\NxR.aluData2[0]~16_combout\ & 
-- \Mux245~0_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100000001000011011100000111001101001100010011110111110001111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux242~0_combout\,
	datab => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datac => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datad => \ALT_INV_Mux245~0_combout\,
	datae => \ALT_INV_Mux244~0_combout\,
	dataf => \ALT_INV_Mux243~0_combout\,
	combout => \ShiftLeft0~16_combout\);

-- Location: FF_X75_Y7_N49
\ShiftLeft0~16_NEW_REG286\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~16_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~16_OTERM287\);

-- Location: LABCELL_X74_Y8_N48
\ShiftLeft0~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~17_combout\ = ( \R.aluData2\(3) & ( \R.aluData2\(2) & ( \ShiftLeft0~0_OTERM263\ ) ) ) # ( !\R.aluData2\(3) & ( \R.aluData2\(2) & ( \ShiftLeft0~10_OTERM211\ ) ) ) # ( \R.aluData2\(3) & ( !\R.aluData2\(2) & ( \ShiftLeft0~5_OTERM203\ ) ) ) # ( 
-- !\R.aluData2\(3) & ( !\R.aluData2\(2) & ( \ShiftLeft0~16_OTERM287\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111000011110000111100110011001100110101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~0_OTERM263\,
	datab => \ALT_INV_ShiftLeft0~10_OTERM211\,
	datac => \ALT_INV_ShiftLeft0~5_OTERM203\,
	datad => \ALT_INV_ShiftLeft0~16_OTERM287\,
	datae => \ALT_INV_R.aluData2\(3),
	dataf => \ALT_INV_R.aluData2\(2),
	combout => \ShiftLeft0~17_combout\);

-- Location: MLABCELL_X84_Y6_N30
\Selector20~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector20~2_combout\ = ( !\R.aluData2\(12) & ( \R.aluOp.ALUOpOr~q\ & ( !\R.aluData1\(12) ) ) ) # ( \R.aluData2\(12) & ( !\R.aluOp.ALUOpOr~q\ & ( (!\R.aluData1\(12) & (!\R.aluOp.ALUOpXor~DUPLICATE_q\)) # (\R.aluData1\(12) & 
-- ((!\R.aluOp.ALUOpAnd~DUPLICATE_q\))) ) ) ) # ( !\R.aluData2\(12) & ( !\R.aluOp.ALUOpOr~q\ & ( (!\R.aluOp.ALUOpXor~DUPLICATE_q\) # (!\R.aluData1\(12)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111101011111010101011111010000011110000111100000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpXor~DUPLICATE_q\,
	datac => \ALT_INV_R.aluData1\(12),
	datad => \ALT_INV_R.aluOp.ALUOpAnd~DUPLICATE_q\,
	datae => \ALT_INV_R.aluData2\(12),
	dataf => \ALT_INV_R.aluOp.ALUOpOr~q\,
	combout => \Selector20~2_combout\);

-- Location: LABCELL_X71_Y7_N54
\Selector20~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector20~0_combout\ = ( \R.aluOp.ALUOpSRA_OTERM363\ & ( (\Mux223~0_combout\ & ((\NxR.aluData2[3]~18_combout\) # (\NxR.aluData2[2]~19_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000101000011110000010100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_NxR.aluData2[2]~19_combout\,
	datac => \ALT_INV_Mux223~0_combout\,
	datad => \ALT_INV_NxR.aluData2[3]~18_combout\,
	dataf => \ALT_INV_R.aluOp.ALUOpSRA_OTERM363\,
	combout => \Selector20~0_combout\);

-- Location: FF_X71_Y7_N55
\Selector20~0_NEW_REG768\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector20~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector20~0_OTERM769\);

-- Location: LABCELL_X73_Y5_N36
\ShiftRight1~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~3_combout\ = ( \NxR.aluData2[0]~16_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( \Mux223~0_combout\ ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( \Mux224~0_combout\ ) ) ) # ( \NxR.aluData2[0]~16_combout\ & ( 
-- !\NxR.aluData2[1]~17_combout\ & ( \Mux225~0_combout\ ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( !\NxR.aluData2[1]~17_combout\ & ( \Mux226~0_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111010101010101010100000000111111110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux225~0_combout\,
	datab => \ALT_INV_Mux223~0_combout\,
	datac => \ALT_INV_Mux226~0_combout\,
	datad => \ALT_INV_Mux224~0_combout\,
	datae => \ALT_INV_NxR.aluData2[0]~16_combout\,
	dataf => \ALT_INV_NxR.aluData2[1]~17_combout\,
	combout => \ShiftRight1~3_combout\);

-- Location: FF_X73_Y5_N37
\ShiftRight1~3_NEW_REG12\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~3_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~3_OTERM13\);

-- Location: MLABCELL_X78_Y4_N39
\Selector20~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector20~1_combout\ = ( \R.aluData2\(4) & ( ((\Selector31~0_OTERM349\ & (\ShiftRight1~3_OTERM13\ & !\ShiftRight0~7_OTERM233DUPLICATE_q\))) # (\Selector20~0_OTERM769\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000001010111010101010101011101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector20~0_OTERM769\,
	datab => \ALT_INV_Selector31~0_OTERM349\,
	datac => \ALT_INV_ShiftRight1~3_OTERM13\,
	datad => \ALT_INV_ShiftRight0~7_OTERM233DUPLICATE_q\,
	dataf => \ALT_INV_R.aluData2\(4),
	combout => \Selector20~1_combout\);

-- Location: LABCELL_X74_Y6_N0
\ShiftRight1~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~0_combout\ = ( \NxR.aluData2[0]~16_combout\ & ( \Mux237~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\) # (\Mux235~0_combout\) ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( \Mux237~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & 
-- ((\Mux238~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux236~0_combout\)) ) ) ) # ( \NxR.aluData2[0]~16_combout\ & ( !\Mux237~0_combout\ & ( (\NxR.aluData2[1]~17_combout\ & \Mux235~0_combout\) ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( 
-- !\Mux237~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((\Mux238~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux236~0_combout\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001101100011011000000000101010100011011000110111010101011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datab => \ALT_INV_Mux236~0_combout\,
	datac => \ALT_INV_Mux238~0_combout\,
	datad => \ALT_INV_Mux235~0_combout\,
	datae => \ALT_INV_NxR.aluData2[0]~16_combout\,
	dataf => \ALT_INV_Mux237~0_combout\,
	combout => \ShiftRight1~0_combout\);

-- Location: FF_X74_Y6_N2
\ShiftRight1~0_NEW_REG256\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~0_OTERM257\);

-- Location: LABCELL_X73_Y8_N33
\ShiftRight1~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~8_combout\ = ( \Mux241~0_combout\ & ( \NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\) # (\Mux239~0_combout\) ) ) ) # ( !\Mux241~0_combout\ & ( \NxR.aluData2[0]~16_combout\ & ( (\NxR.aluData2[1]~17_combout\ & 
-- \Mux239~0_combout\) ) ) ) # ( \Mux241~0_combout\ & ( !\NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (\Mux242~0_combout\)) # (\NxR.aluData2[1]~17_combout\ & ((\Mux240~0_combout\))) ) ) ) # ( !\Mux241~0_combout\ & ( 
-- !\NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (\Mux242~0_combout\)) # (\NxR.aluData2[1]~17_combout\ & ((\Mux240~0_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010011100100111001001110010011100000000010101011010101011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datab => \ALT_INV_Mux242~0_combout\,
	datac => \ALT_INV_Mux240~0_combout\,
	datad => \ALT_INV_Mux239~0_combout\,
	datae => \ALT_INV_Mux241~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[0]~16_combout\,
	combout => \ShiftRight1~8_combout\);

-- Location: FF_X73_Y8_N34
\ShiftRight1~8_NEW_REG260\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~8_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~8_OTERM261\);

-- Location: LABCELL_X74_Y3_N42
\ShiftRight1~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~1_combout\ = ( \Mux234~0_combout\ & ( \NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((\Mux233~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux231~0_combout\)) ) ) ) # ( !\Mux234~0_combout\ & ( 
-- \NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((\Mux233~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux231~0_combout\)) ) ) ) # ( \Mux234~0_combout\ & ( !\NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\) # 
-- (\Mux232~0_combout\) ) ) ) # ( !\Mux234~0_combout\ & ( !\NxR.aluData2[0]~16_combout\ & ( (\Mux232~0_combout\ & \NxR.aluData2[1]~17_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010101111111110101010100001111001100110000111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux232~0_combout\,
	datab => \ALT_INV_Mux231~0_combout\,
	datac => \ALT_INV_Mux233~0_combout\,
	datad => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datae => \ALT_INV_Mux234~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[0]~16_combout\,
	combout => \ShiftRight1~1_combout\);

-- Location: FF_X74_Y3_N43
\ShiftRight1~1_NEW_REG32\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~1_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~1_OTERM33\);

-- Location: LABCELL_X74_Y5_N45
\ShiftRight1~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~2_combout\ = ( \Mux230~0_combout\ & ( \NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((\Mux229~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux227~0_combout\)) ) ) ) # ( !\Mux230~0_combout\ & ( 
-- \NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((\Mux229~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux227~0_combout\)) ) ) ) # ( \Mux230~0_combout\ & ( !\NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\) # 
-- (\Mux228~0_combout\) ) ) ) # ( !\Mux230~0_combout\ & ( !\NxR.aluData2[0]~16_combout\ & ( (\NxR.aluData2[1]~17_combout\ & \Mux228~0_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110011110011001111111100011101000111010001110100011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux227~0_combout\,
	datab => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datac => \ALT_INV_Mux229~0_combout\,
	datad => \ALT_INV_Mux228~0_combout\,
	datae => \ALT_INV_Mux230~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[0]~16_combout\,
	combout => \ShiftRight1~2_combout\);

-- Location: FF_X74_Y5_N46
\ShiftRight1~2_NEW_REG48\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~2_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~2_OTERM49\);

-- Location: LABCELL_X75_Y8_N24
\ShiftRight1~51\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~51_combout\ = ( \R.aluData2\(3) & ( \R.aluData2\(2) & ( \ShiftRight1~2_OTERM49\ ) ) ) # ( !\R.aluData2\(3) & ( \R.aluData2\(2) & ( \ShiftRight1~0_OTERM257\ ) ) ) # ( \R.aluData2\(3) & ( !\R.aluData2\(2) & ( \ShiftRight1~1_OTERM33\ ) ) ) # ( 
-- !\R.aluData2\(3) & ( !\R.aluData2\(2) & ( \ShiftRight1~8_OTERM261\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110011000011110000111101010101010101010000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~0_OTERM257\,
	datab => \ALT_INV_ShiftRight1~8_OTERM261\,
	datac => \ALT_INV_ShiftRight1~1_OTERM33\,
	datad => \ALT_INV_ShiftRight1~2_OTERM49\,
	datae => \ALT_INV_R.aluData2\(3),
	dataf => \ALT_INV_R.aluData2\(2),
	combout => \ShiftRight1~51_combout\);

-- Location: LABCELL_X81_Y4_N18
\Selector20~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector20~3_combout\ = ( !\Selector20~1_combout\ & ( \ShiftRight1~51_combout\ & ( (\Selector20~2_combout\ & (!\Selector31~5_OTERM599\ & ((!\Selector27~0_OTERM385\) # (!\ShiftLeft0~17_combout\)))) ) ) ) # ( !\Selector20~1_combout\ & ( 
-- !\ShiftRight1~51_combout\ & ( (\Selector20~2_combout\ & ((!\Selector27~0_OTERM385\) # (!\ShiftLeft0~17_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111000001110000000000000000000001110000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector27~0_OTERM385\,
	datab => \ALT_INV_ShiftLeft0~17_combout\,
	datac => \ALT_INV_Selector20~2_combout\,
	datad => \ALT_INV_Selector31~5_OTERM599\,
	datae => \ALT_INV_Selector20~1_combout\,
	dataf => \ALT_INV_ShiftRight1~51_combout\,
	combout => \Selector20~3_combout\);

-- Location: LABCELL_X74_Y3_N36
\ShiftRight1~31\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~31_combout\ = ( \NxR.aluData2[0]~16_combout\ & ( \Mux229~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((\Mux230~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux228~0_combout\)) ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( 
-- \Mux229~0_combout\ & ( (\NxR.aluData2[1]~17_combout\) # (\Mux231~0_combout\) ) ) ) # ( \NxR.aluData2[0]~16_combout\ & ( !\Mux229~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((\Mux230~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & 
-- (\Mux228~0_combout\)) ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( !\Mux229~0_combout\ & ( (\Mux231~0_combout\ & !\NxR.aluData2[1]~17_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010100000000000011110011001101010101111111110000111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux231~0_combout\,
	datab => \ALT_INV_Mux228~0_combout\,
	datac => \ALT_INV_Mux230~0_combout\,
	datad => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datae => \ALT_INV_NxR.aluData2[0]~16_combout\,
	dataf => \ALT_INV_Mux229~0_combout\,
	combout => \ShiftRight1~31_combout\);

-- Location: FF_X74_Y3_N37
\ShiftRight1~31_NEW_REG44\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~31_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~31_OTERM45\);

-- Location: LABCELL_X80_Y7_N33
\Selector25~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector25~2_combout\ = ( \ShiftRight1~31_OTERM45\ & ( \R.aluData2\(3) & ( (\ShiftRight0~4_OTERM31\ & (\Selector31~7_OTERM383\ & !\R.aluData2\(2))) ) ) ) # ( !\ShiftRight1~31_OTERM45\ & ( \R.aluData2\(3) & ( (\ShiftRight0~4_OTERM31\ & 
-- (\Selector31~7_OTERM383\ & !\R.aluData2\(2))) ) ) ) # ( \ShiftRight1~31_OTERM45\ & ( !\R.aluData2\(3) & ( (\Selector31~7_OTERM383\ & ((!\R.aluData2\(2)) # (\ShiftRight1~32_OTERM21\))) ) ) ) # ( !\ShiftRight1~31_OTERM45\ & ( !\R.aluData2\(3) & ( 
-- (\ShiftRight1~32_OTERM21\ & (\Selector31~7_OTERM383\ & \R.aluData2\(2))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000011000011110000001100000101000000000000010100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight0~4_OTERM31\,
	datab => \ALT_INV_ShiftRight1~32_OTERM21\,
	datac => \ALT_INV_Selector31~7_OTERM383\,
	datad => \ALT_INV_R.aluData2\(2),
	datae => \ALT_INV_ShiftRight1~31_OTERM45\,
	dataf => \ALT_INV_R.aluData2\(3),
	combout => \Selector25~2_combout\);

-- Location: LABCELL_X74_Y5_N30
\ShiftRight1~30\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~30_combout\ = ( \NxR.aluData2[1]~17_combout\ & ( \Mux232~0_combout\ & ( (\NxR.aluData2[0]~16_combout\) # (\Mux233~0_combout\) ) ) ) # ( !\NxR.aluData2[1]~17_combout\ & ( \Mux232~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & 
-- (\Mux235~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & ((\Mux234~0_combout\))) ) ) ) # ( \NxR.aluData2[1]~17_combout\ & ( !\Mux232~0_combout\ & ( (\Mux233~0_combout\ & !\NxR.aluData2[0]~16_combout\) ) ) ) # ( !\NxR.aluData2[1]~17_combout\ & ( 
-- !\Mux232~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (\Mux235~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & ((\Mux234~0_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011000000111111010100000101000000110000001111110101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux233~0_combout\,
	datab => \ALT_INV_Mux235~0_combout\,
	datac => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datad => \ALT_INV_Mux234~0_combout\,
	datae => \ALT_INV_NxR.aluData2[1]~17_combout\,
	dataf => \ALT_INV_Mux232~0_combout\,
	combout => \ShiftRight1~30_combout\);

-- Location: FF_X74_Y5_N31
\ShiftRight1~30_NEW_REG38\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~30_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~30_OTERM39\);

-- Location: LABCELL_X73_Y6_N12
\ShiftRight1~37\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~37_combout\ = ( \Mux236~0_combout\ & ( \Mux239~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (((!\NxR.aluData2[1]~17_combout\)) # (\Mux237~0_combout\))) # (\NxR.aluData2[0]~16_combout\ & (((\NxR.aluData2[1]~17_combout\) # 
-- (\Mux238~0_combout\)))) ) ) ) # ( !\Mux236~0_combout\ & ( \Mux239~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (((!\NxR.aluData2[1]~17_combout\)) # (\Mux237~0_combout\))) # (\NxR.aluData2[0]~16_combout\ & (((\Mux238~0_combout\ & 
-- !\NxR.aluData2[1]~17_combout\)))) ) ) ) # ( \Mux236~0_combout\ & ( !\Mux239~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (\Mux237~0_combout\ & ((\NxR.aluData2[1]~17_combout\)))) # (\NxR.aluData2[0]~16_combout\ & (((\NxR.aluData2[1]~17_combout\) # 
-- (\Mux238~0_combout\)))) ) ) ) # ( !\Mux236~0_combout\ & ( !\Mux239~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (\Mux237~0_combout\ & ((\NxR.aluData2[1]~17_combout\)))) # (\NxR.aluData2[0]~16_combout\ & (((\Mux238~0_combout\ & 
-- !\NxR.aluData2[1]~17_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001101000100000000110111011111001111010001001100111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux237~0_combout\,
	datab => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datac => \ALT_INV_Mux238~0_combout\,
	datad => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datae => \ALT_INV_Mux236~0_combout\,
	dataf => \ALT_INV_Mux239~0_combout\,
	combout => \ShiftRight1~37_combout\);

-- Location: FF_X73_Y6_N13
\ShiftRight1~37_NEW_REG282\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~37_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~37_OTERM283\);

-- Location: LABCELL_X75_Y7_N42
\ShiftRight1~35\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~35_combout\ = ( \Mux244~0_combout\ & ( \Mux247~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (((!\NxR.aluData2[1]~17_combout\) # (\Mux245~0_combout\)))) # (\NxR.aluData2[0]~16_combout\ & (((\NxR.aluData2[1]~17_combout\)) # 
-- (\Mux246~0_combout\))) ) ) ) # ( !\Mux244~0_combout\ & ( \Mux247~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (((!\NxR.aluData2[1]~17_combout\) # (\Mux245~0_combout\)))) # (\NxR.aluData2[0]~16_combout\ & (\Mux246~0_combout\ & 
-- ((!\NxR.aluData2[1]~17_combout\)))) ) ) ) # ( \Mux244~0_combout\ & ( !\Mux247~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (((\Mux245~0_combout\ & \NxR.aluData2[1]~17_combout\)))) # (\NxR.aluData2[0]~16_combout\ & (((\NxR.aluData2[1]~17_combout\)) # 
-- (\Mux246~0_combout\))) ) ) ) # ( !\Mux244~0_combout\ & ( !\Mux247~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (((\Mux245~0_combout\ & \NxR.aluData2[1]~17_combout\)))) # (\NxR.aluData2[0]~16_combout\ & (\Mux246~0_combout\ & 
-- ((!\NxR.aluData2[1]~17_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100110000000001010011111111110101001100001111010100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux246~0_combout\,
	datab => \ALT_INV_Mux245~0_combout\,
	datac => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datad => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datae => \ALT_INV_Mux244~0_combout\,
	dataf => \ALT_INV_Mux247~0_combout\,
	combout => \ShiftRight1~35_combout\);

-- Location: FF_X75_Y7_N43
\ShiftRight1~35_NEW_REG278\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~35_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~35_OTERM279\);

-- Location: LABCELL_X77_Y7_N48
\ShiftRight1~45\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~45_combout\ = ( \ShiftRight1~35_OTERM279\ & ( \ShiftRight1~36_OTERM281\ & ( (!\R.aluData2\(3)) # ((!\R.aluData2\(2) & ((\ShiftRight1~37_OTERM283\))) # (\R.aluData2\(2) & (\ShiftRight1~30_OTERM39\))) ) ) ) # ( !\ShiftRight1~35_OTERM279\ & ( 
-- \ShiftRight1~36_OTERM281\ & ( (!\R.aluData2\(2) & (((\ShiftRight1~37_OTERM283\ & \R.aluData2\(3))))) # (\R.aluData2\(2) & (((!\R.aluData2\(3))) # (\ShiftRight1~30_OTERM39\))) ) ) ) # ( \ShiftRight1~35_OTERM279\ & ( !\ShiftRight1~36_OTERM281\ & ( 
-- (!\R.aluData2\(2) & (((!\R.aluData2\(3)) # (\ShiftRight1~37_OTERM283\)))) # (\R.aluData2\(2) & (\ShiftRight1~30_OTERM39\ & ((\R.aluData2\(3))))) ) ) ) # ( !\ShiftRight1~35_OTERM279\ & ( !\ShiftRight1~36_OTERM281\ & ( (\R.aluData2\(3) & ((!\R.aluData2\(2) 
-- & ((\ShiftRight1~37_OTERM283\))) # (\R.aluData2\(2) & (\ShiftRight1~30_OTERM39\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000011101110011000001110100110011000111011111111100011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~30_OTERM39\,
	datab => \ALT_INV_R.aluData2\(2),
	datac => \ALT_INV_ShiftRight1~37_OTERM283\,
	datad => \ALT_INV_R.aluData2\(3),
	datae => \ALT_INV_ShiftRight1~35_OTERM279\,
	dataf => \ALT_INV_ShiftRight1~36_OTERM281\,
	combout => \ShiftRight1~45_combout\);

-- Location: LABCELL_X74_Y7_N30
\Selector25~3_RTM0799\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector25~3_RTM0799_combout\ = ( \NxR.aluData2[7]~14_combout\ & ( ((!\Mux247~0_combout\ & (\R.aluOp.ALUOpXor_OTERM355\)) # (\Mux247~0_combout\ & ((\R.aluOp.ALUOpAnd_OTERM357\)))) # (\R.aluOp.ALUOpOr_OTERM353\) ) ) # ( !\NxR.aluData2[7]~14_combout\ & ( 
-- (\Mux247~0_combout\ & ((\R.aluOp.ALUOpXor_OTERM355\) # (\R.aluOp.ALUOpOr_OTERM353\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001110111000000000111011101110111010111110111011101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpOr_OTERM353\,
	datab => \ALT_INV_R.aluOp.ALUOpXor_OTERM355\,
	datac => \ALT_INV_R.aluOp.ALUOpAnd_OTERM357\,
	datad => \ALT_INV_Mux247~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[7]~14_combout\,
	combout => \Selector25~3_RTM0799_combout\);

-- Location: FF_X74_Y7_N32
\Selector25~3_NEW_REG796\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector25~3_RTM0799_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector25~3_OTERM797\);

-- Location: LABCELL_X80_Y7_N51
\Selector25~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector25~4_combout\ = ( \ShiftLeft0~3_OTERM223\ & ( \R.aluData2\(3) & ( !\Selector25~3_OTERM797\ ) ) ) # ( !\ShiftLeft0~3_OTERM223\ & ( \R.aluData2\(3) & ( !\Selector25~3_OTERM797\ ) ) ) # ( \ShiftLeft0~3_OTERM223\ & ( !\R.aluData2\(3) & ( 
-- (!\Selector25~3_OTERM797\ & ((!\Selector27~0_OTERM385\) # ((!\R.aluData2\(2) & !\ShiftLeft0~9_OTERM461\)))) ) ) ) # ( !\ShiftLeft0~3_OTERM223\ & ( !\R.aluData2\(3) & ( (!\Selector25~3_OTERM797\ & (((!\ShiftLeft0~9_OTERM461\) # (!\Selector27~0_OTERM385\)) 
-- # (\R.aluData2\(2)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010101010100010101010101000000010101010101010101010101010101010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector25~3_OTERM797\,
	datab => \ALT_INV_R.aluData2\(2),
	datac => \ALT_INV_ShiftLeft0~9_OTERM461\,
	datad => \ALT_INV_Selector27~0_OTERM385\,
	datae => \ALT_INV_ShiftLeft0~3_OTERM223\,
	dataf => \ALT_INV_R.aluData2\(3),
	combout => \Selector25~4_combout\);

-- Location: LABCELL_X83_Y5_N18
\Selector25~6_RESYN1116\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector25~6_RESYN1116_BDD1117\ = ( \ShiftRight1~45_combout\ & ( \Selector25~4_combout\ & ( (\Selector25~2_combout\) # (\Selector31~5_OTERM599\) ) ) ) # ( !\ShiftRight1~45_combout\ & ( \Selector25~4_combout\ & ( \Selector25~2_combout\ ) ) ) # ( 
-- \ShiftRight1~45_combout\ & ( !\Selector25~4_combout\ ) ) # ( !\ShiftRight1~45_combout\ & ( !\Selector25~4_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111111111111111111100001111000011110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Selector31~5_OTERM599\,
	datac => \ALT_INV_Selector25~2_combout\,
	datae => \ALT_INV_ShiftRight1~45_combout\,
	dataf => \ALT_INV_Selector25~4_combout\,
	combout => \Selector25~6_RESYN1116_BDD1117\);

-- Location: LABCELL_X77_Y9_N51
\Selector25~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector25~1_combout\ = ( \ShiftRight1~31_OTERM45\ & ( \ShiftRight1~32_OTERM21\ & ( (\Selector31~6_OTERM381\ & ((!\R.aluData2\(3)) # (\R.aluData1\(31)))) ) ) ) # ( !\ShiftRight1~31_OTERM45\ & ( \ShiftRight1~32_OTERM21\ & ( (\Selector31~6_OTERM381\ & 
-- ((!\R.aluData2\(3) & ((\R.aluData2\(2)))) # (\R.aluData2\(3) & (\R.aluData1\(31))))) ) ) ) # ( \ShiftRight1~31_OTERM45\ & ( !\ShiftRight1~32_OTERM21\ & ( (\Selector31~6_OTERM381\ & ((!\R.aluData2\(3) & ((!\R.aluData2\(2)))) # (\R.aluData2\(3) & 
-- (\R.aluData1\(31))))) ) ) ) # ( !\ShiftRight1~31_OTERM45\ & ( !\ShiftRight1~32_OTERM21\ & ( (\R.aluData1\(31) & (\Selector31~6_OTERM381\ & \R.aluData2\(3))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000101000011000000010100000011000001010000111100000101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData1\(31),
	datab => \ALT_INV_R.aluData2\(2),
	datac => \ALT_INV_Selector31~6_OTERM381\,
	datad => \ALT_INV_R.aluData2\(3),
	datae => \ALT_INV_ShiftRight1~31_OTERM45\,
	dataf => \ALT_INV_ShiftRight1~32_OTERM21\,
	combout => \Selector25~1_combout\);

-- Location: LABCELL_X83_Y5_N54
\Selector25~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector25~6_combout\ = ( \R.aluOp.ALUOpSub~q\ & ( \Add2~29_sumout\ ) ) # ( !\R.aluOp.ALUOpSub~q\ & ( \Add2~29_sumout\ & ( (((\R.aluOp.ALUOpAdd~q\ & \Add1~29_sumout\)) # (\Selector25~1_combout\)) # (\Selector25~6_RESYN1116_BDD1117\) ) ) ) # ( 
-- \R.aluOp.ALUOpSub~q\ & ( !\Add2~29_sumout\ & ( (((\R.aluOp.ALUOpAdd~q\ & \Add1~29_sumout\)) # (\Selector25~1_combout\)) # (\Selector25~6_RESYN1116_BDD1117\) ) ) ) # ( !\R.aluOp.ALUOpSub~q\ & ( !\Add2~29_sumout\ & ( (((\R.aluOp.ALUOpAdd~q\ & 
-- \Add1~29_sumout\)) # (\Selector25~1_combout\)) # (\Selector25~6_RESYN1116_BDD1117\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001111111111111000111111111111100011111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datab => \ALT_INV_Add1~29_sumout\,
	datac => \ALT_INV_Selector25~6_RESYN1116_BDD1117\,
	datad => \ALT_INV_Selector25~1_combout\,
	datae => \ALT_INV_R.aluOp.ALUOpSub~q\,
	dataf => \ALT_INV_Add2~29_sumout\,
	combout => \Selector25~6_combout\);

-- Location: MLABCELL_X78_Y6_N36
\Add1~49\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~49_sumout\ = SUM(( \R.aluData2\(12) ) + ( \R.aluData1\(12) ) + ( \Add1~46\ ))
-- \Add1~50\ = CARRY(( \R.aluData2\(12) ) + ( \R.aluData1\(12) ) + ( \Add1~46\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluData2\(12),
	datac => \ALT_INV_R.aluData1\(12),
	cin => \Add1~46\,
	sumout => \Add1~49_sumout\,
	cout => \Add1~50\);

-- Location: LABCELL_X81_Y4_N45
\Selector20~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector20~6_combout\ = ( \R.aluOp.ALUOpSub~q\ & ( (!\Selector20~3_combout\) # (((\Add1~49_sumout\ & \R.aluOp.ALUOpAdd~q\)) # (\Add2~49_sumout\)) ) ) # ( !\R.aluOp.ALUOpSub~q\ & ( (!\Selector20~3_combout\) # ((\Add1~49_sumout\ & \R.aluOp.ALUOpAdd~q\)) ) 
-- )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010101010101111101010101010111110111011101111111011101110111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector20~3_combout\,
	datab => \ALT_INV_Add2~49_sumout\,
	datac => \ALT_INV_Add1~49_sumout\,
	datad => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	dataf => \ALT_INV_R.aluOp.ALUOpSub~q\,
	combout => \Selector20~6_combout\);

-- Location: FF_X81_Y4_N47
\R.aluRes[12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector20~6_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(12));

-- Location: FF_X83_Y5_N56
\R.aluRes[7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector25~6_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(7));

-- Location: LABCELL_X81_Y4_N30
\Equal3~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \Equal3~10_combout\ = ( \Add1~49_sumout\ & ( \R.aluCalc~q\ & ( !\R.aluOp.ALUOpAdd~q\ ) ) ) # ( !\Add1~49_sumout\ & ( \R.aluCalc~q\ ) ) # ( \Add1~49_sumout\ & ( !\R.aluCalc~q\ & ( (!\R.aluRes\(12) & !\R.aluRes\(7)) ) ) ) # ( !\Add1~49_sumout\ & ( 
-- !\R.aluCalc~q\ & ( (!\R.aluRes\(12) & !\R.aluRes\(7)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1100000011000000110000001100000011111111111111111111111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluRes\(12),
	datac => \ALT_INV_R.aluRes\(7),
	datad => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datae => \ALT_INV_Add1~49_sumout\,
	dataf => \ALT_INV_R.aluCalc~q\,
	combout => \Equal3~10_combout\);

-- Location: LABCELL_X81_Y4_N48
\Equal3~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Equal3~3_combout\ = ( \Add2~49_sumout\ & ( \R.aluOp.ALUOpSub~q\ & ( (!\R.aluCalc~q\ & \Equal3~10_combout\) ) ) ) # ( !\Add2~49_sumout\ & ( \R.aluOp.ALUOpSub~q\ & ( (\Equal3~10_combout\ & ((!\R.aluCalc~q\) # ((\Selector20~3_combout\ & 
-- !\Selector25~6_combout\)))) ) ) ) # ( \Add2~49_sumout\ & ( !\R.aluOp.ALUOpSub~q\ & ( (\Equal3~10_combout\ & ((!\R.aluCalc~q\) # ((\Selector20~3_combout\ & !\Selector25~6_combout\)))) ) ) ) # ( !\Add2~49_sumout\ & ( !\R.aluOp.ALUOpSub~q\ & ( 
-- (\Equal3~10_combout\ & ((!\R.aluCalc~q\) # ((\Selector20~3_combout\ & !\Selector25~6_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011110100000000001111010000000000111101000000000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector20~3_combout\,
	datab => \ALT_INV_Selector25~6_combout\,
	datac => \ALT_INV_R.aluCalc~q\,
	datad => \ALT_INV_Equal3~10_combout\,
	datae => \ALT_INV_Add2~49_sumout\,
	dataf => \ALT_INV_R.aluOp.ALUOpSub~q\,
	combout => \Equal3~3_combout\);

-- Location: FF_X81_Y4_N49
\R.statusReg[0]_OTERM9_NEW_REG468\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Equal3~3_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.statusReg[0]_OTERM9_OTERM469\);

-- Location: LABCELL_X77_Y8_N15
\LessThan1~31\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~31_combout\ = ( \R.aluData1\(22) & ( !\R.aluData2\(22) ) ) # ( !\R.aluData1\(22) & ( \R.aluData2\(22) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111000000001111111111111111000000001111111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \ALT_INV_R.aluData2\(22),
	dataf => \ALT_INV_R.aluData1\(22),
	combout => \LessThan1~31_combout\);

-- Location: LABCELL_X77_Y8_N18
\Selector10~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector10~2_combout\ = ( \ShiftLeft0~8_OTERM207\ & ( (!\R.aluData2\(3) & (\Selector12~2_OTERM395\ & ((!\R.aluData2\(2)) # (\ShiftLeft0~2_OTERM221\)))) ) ) # ( !\ShiftLeft0~8_OTERM207\ & ( (!\R.aluData2\(3) & (\R.aluData2\(2) & (\ShiftLeft0~2_OTERM221\ & 
-- \Selector12~2_OTERM395\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000010000000000000001000000000100010100000000010001010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(3),
	datab => \ALT_INV_R.aluData2\(2),
	datac => \ALT_INV_ShiftLeft0~2_OTERM221\,
	datad => \ALT_INV_Selector12~2_OTERM395\,
	dataf => \ALT_INV_ShiftLeft0~8_OTERM207\,
	combout => \Selector10~2_combout\);

-- Location: LABCELL_X77_Y8_N33
\Selector10~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector10~3_combout\ = ( \R.aluOp.ALUOpOr~q\ & ( (\R.aluData2\(22)) # (\R.aluData1\(22)) ) ) # ( !\R.aluOp.ALUOpOr~q\ & ( (\R.aluOp.ALUOpAnd~DUPLICATE_q\ & (\R.aluData1\(22) & \R.aluData2\(22))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000101000000000000010100001111111111110000111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpAnd~DUPLICATE_q\,
	datac => \ALT_INV_R.aluData1\(22),
	datad => \ALT_INV_R.aluData2\(22),
	dataf => \ALT_INV_R.aluOp.ALUOpOr~q\,
	combout => \Selector10~3_combout\);

-- Location: LABCELL_X77_Y8_N24
\Selector10~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector10~4_combout\ = ( !\Selector10~3_combout\ & ( (!\Selector17~0_OTERM391\ & (!\Selector10~2_combout\ & ((!\LessThan1~31_combout\) # (!\R.aluOp.ALUOpXor~DUPLICATE_q\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010000010000000101000001000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector17~0_OTERM391\,
	datab => \ALT_INV_LessThan1~31_combout\,
	datac => \ALT_INV_Selector10~2_combout\,
	datad => \ALT_INV_R.aluOp.ALUOpXor~DUPLICATE_q\,
	dataf => \ALT_INV_Selector10~3_combout\,
	combout => \Selector10~4_combout\);

-- Location: LABCELL_X74_Y6_N24
\ShiftLeft0~20\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~20_combout\ = ( \Mux243~0_combout\ & ( \NxR.aluData2[0]~16_combout\ & ( (\NxR.aluData2[1]~17_combout\) # (\Mux241~0_combout\) ) ) ) # ( !\Mux243~0_combout\ & ( \NxR.aluData2[0]~16_combout\ & ( (\Mux241~0_combout\ & 
-- !\NxR.aluData2[1]~17_combout\) ) ) ) # ( \Mux243~0_combout\ & ( !\NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (\Mux240~0_combout\)) # (\NxR.aluData2[1]~17_combout\ & ((\Mux242~0_combout\))) ) ) ) # ( !\Mux243~0_combout\ & ( 
-- !\NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (\Mux240~0_combout\)) # (\NxR.aluData2[1]~17_combout\ & ((\Mux242~0_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010100001111010101010000111100110011000000000011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux240~0_combout\,
	datab => \ALT_INV_Mux241~0_combout\,
	datac => \ALT_INV_Mux242~0_combout\,
	datad => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datae => \ALT_INV_Mux243~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[0]~16_combout\,
	combout => \ShiftLeft0~20_combout\);

-- Location: FF_X74_Y6_N25
\ShiftLeft0~20_NEW_REG290\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~20_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~20_OTERM291\);

-- Location: LABCELL_X75_Y7_N15
\ShiftLeft0~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~13_combout\ = ( \Mux244~0_combout\ & ( \Mux247~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((!\NxR.aluData2[0]~16_combout\) # (\Mux245~0_combout\)))) # (\NxR.aluData2[1]~17_combout\ & (((\NxR.aluData2[0]~16_combout\)) # 
-- (\Mux246~0_combout\))) ) ) ) # ( !\Mux244~0_combout\ & ( \Mux247~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((\Mux245~0_combout\ & \NxR.aluData2[0]~16_combout\)))) # (\NxR.aluData2[1]~17_combout\ & (((\NxR.aluData2[0]~16_combout\)) # 
-- (\Mux246~0_combout\))) ) ) ) # ( \Mux244~0_combout\ & ( !\Mux247~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((!\NxR.aluData2[0]~16_combout\) # (\Mux245~0_combout\)))) # (\NxR.aluData2[1]~17_combout\ & (\Mux246~0_combout\ & 
-- ((!\NxR.aluData2[0]~16_combout\)))) ) ) ) # ( !\Mux244~0_combout\ & ( !\Mux247~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((\Mux245~0_combout\ & \NxR.aluData2[0]~16_combout\)))) # (\NxR.aluData2[1]~17_combout\ & (\Mux246~0_combout\ & 
-- ((!\NxR.aluData2[0]~16_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100110000111101010011000000000101001111111111010100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux246~0_combout\,
	datab => \ALT_INV_Mux245~0_combout\,
	datac => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datad => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datae => \ALT_INV_Mux244~0_combout\,
	dataf => \ALT_INV_Mux247~0_combout\,
	combout => \ShiftLeft0~13_combout\);

-- Location: FF_X75_Y7_N16
\ShiftLeft0~13_NEW_REG284\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~13_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~13_OTERM285\);

-- Location: LABCELL_X73_Y6_N24
\ShiftLeft0~28\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~28_combout\ = ( \Mux236~0_combout\ & ( \Mux239~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (((!\NxR.aluData2[1]~17_combout\) # (\Mux238~0_combout\)))) # (\NxR.aluData2[0]~16_combout\ & (((\NxR.aluData2[1]~17_combout\)) # 
-- (\Mux237~0_combout\))) ) ) ) # ( !\Mux236~0_combout\ & ( \Mux239~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (((\Mux238~0_combout\ & \NxR.aluData2[1]~17_combout\)))) # (\NxR.aluData2[0]~16_combout\ & (((\NxR.aluData2[1]~17_combout\)) # 
-- (\Mux237~0_combout\))) ) ) ) # ( \Mux236~0_combout\ & ( !\Mux239~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (((!\NxR.aluData2[1]~17_combout\) # (\Mux238~0_combout\)))) # (\NxR.aluData2[0]~16_combout\ & (\Mux237~0_combout\ & 
-- ((!\NxR.aluData2[1]~17_combout\)))) ) ) ) # ( !\Mux236~0_combout\ & ( !\Mux239~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (((\Mux238~0_combout\ & \NxR.aluData2[1]~17_combout\)))) # (\NxR.aluData2[0]~16_combout\ & (\Mux237~0_combout\ & 
-- ((!\NxR.aluData2[1]~17_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100001100110111010000110000010001001111111101110100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux237~0_combout\,
	datab => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datac => \ALT_INV_Mux238~0_combout\,
	datad => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datae => \ALT_INV_Mux236~0_combout\,
	dataf => \ALT_INV_Mux239~0_combout\,
	combout => \ShiftLeft0~28_combout\);

-- Location: FF_X73_Y6_N25
\ShiftLeft0~28_NEW_REG294\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~28_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~28_OTERM295\);

-- Location: LABCELL_X75_Y3_N6
\ShiftLeft0~37\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~37_combout\ = ( \ShiftLeft0~28_OTERM295\ & ( \ShiftLeft0~36_OTERM603\ & ( (!\R.aluData2\(3)) # ((!\R.aluData2\(2) & (\ShiftLeft0~20_OTERM291\)) # (\R.aluData2\(2) & ((\ShiftLeft0~13_OTERM285\)))) ) ) ) # ( !\ShiftLeft0~28_OTERM295\ & ( 
-- \ShiftLeft0~36_OTERM603\ & ( (!\R.aluData2\(2) & (((!\R.aluData2\(3))) # (\ShiftLeft0~20_OTERM291\))) # (\R.aluData2\(2) & (((\ShiftLeft0~13_OTERM285\ & \R.aluData2\(3))))) ) ) ) # ( \ShiftLeft0~28_OTERM295\ & ( !\ShiftLeft0~36_OTERM603\ & ( 
-- (!\R.aluData2\(2) & (\ShiftLeft0~20_OTERM291\ & ((\R.aluData2\(3))))) # (\R.aluData2\(2) & (((!\R.aluData2\(3)) # (\ShiftLeft0~13_OTERM285\)))) ) ) ) # ( !\ShiftLeft0~28_OTERM295\ & ( !\ShiftLeft0~36_OTERM603\ & ( (\R.aluData2\(3) & ((!\R.aluData2\(2) & 
-- (\ShiftLeft0~20_OTERM291\)) # (\R.aluData2\(2) & ((\ShiftLeft0~13_OTERM285\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001000111001100110100011111001100010001111111111101000111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~20_OTERM291\,
	datab => \ALT_INV_R.aluData2\(2),
	datac => \ALT_INV_ShiftLeft0~13_OTERM285\,
	datad => \ALT_INV_R.aluData2\(3),
	datae => \ALT_INV_ShiftLeft0~28_OTERM295\,
	dataf => \ALT_INV_ShiftLeft0~36_OTERM603\,
	combout => \ShiftLeft0~37_combout\);

-- Location: LABCELL_X71_Y6_N24
\ShiftRight0~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight0~2_combout\ = ( \NxR.aluData2[0]~16_combout\ & ( \Mux224~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & \Mux223~0_combout\) ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( \Mux224~0_combout\ & ( !\NxR.aluData2[1]~17_combout\ ) ) ) # ( 
-- \NxR.aluData2[0]~16_combout\ & ( !\Mux224~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & \Mux223~0_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000001111000011110000111100000000000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datad => \ALT_INV_Mux223~0_combout\,
	datae => \ALT_INV_NxR.aluData2[0]~16_combout\,
	dataf => \ALT_INV_Mux224~0_combout\,
	combout => \ShiftRight0~2_combout\);

-- Location: FF_X71_Y6_N25
\ShiftRight0~2_NEW_REG24\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight0~2_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight0~2_OTERM25\);

-- Location: MLABCELL_X82_Y6_N30
\Selector10~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector10~0_combout\ = ( \R.aluData2\(2) & ( \ShiftRight1~27_OTERM19\ & ( (\R.aluOp.ALUOpSRL~q\ & !\R.aluData2\(3)) ) ) ) # ( !\R.aluData2\(2) & ( \ShiftRight1~27_OTERM19\ & ( (\R.aluOp.ALUOpSRL~q\ & ((!\R.aluData2\(3) & (\ShiftRight1~26_OTERM37\)) # 
-- (\R.aluData2\(3) & ((\ShiftRight0~2_OTERM25\))))) ) ) ) # ( !\R.aluData2\(2) & ( !\ShiftRight1~27_OTERM19\ & ( (\R.aluOp.ALUOpSRL~q\ & ((!\R.aluData2\(3) & (\ShiftRight1~26_OTERM37\)) # (\R.aluData2\(3) & ((\ShiftRight0~2_OTERM25\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000011000000000000000000000101000000110000111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~26_OTERM37\,
	datab => \ALT_INV_ShiftRight0~2_OTERM25\,
	datac => \ALT_INV_R.aluOp.ALUOpSRL~q\,
	datad => \ALT_INV_R.aluData2\(3),
	datae => \ALT_INV_R.aluData2\(2),
	dataf => \ALT_INV_ShiftRight1~27_OTERM19\,
	combout => \Selector10~0_combout\);

-- Location: LABCELL_X77_Y2_N30
\Selector10~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector10~1_combout\ = ( !\R.aluData2\(4) & ( \Selector10~0_combout\ ) ) # ( !\R.aluData2\(4) & ( !\Selector10~0_combout\ & ( (!\ShiftLeft0~37_combout\ & (\R.aluOp.ALUOpSRA~q\ & (\ShiftRight1~43_combout\))) # (\ShiftLeft0~37_combout\ & 
-- (((\R.aluOp.ALUOpSRA~q\ & \ShiftRight1~43_combout\)) # (\R.aluOp.ALUOpSLL~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001101010111000000000000000011111111111111110000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~37_combout\,
	datab => \ALT_INV_R.aluOp.ALUOpSRA~q\,
	datac => \ALT_INV_ShiftRight1~43_combout\,
	datad => \ALT_INV_R.aluOp.ALUOpSLL~q\,
	datae => \ALT_INV_R.aluData2\(4),
	dataf => \ALT_INV_Selector10~0_combout\,
	combout => \Selector10~1_combout\);

-- Location: LABCELL_X77_Y2_N48
\Selector10~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector10~5_combout\ = ( \R.aluOp.ALUOpAdd~q\ & ( \Add1~89_sumout\ ) ) # ( !\R.aluOp.ALUOpAdd~q\ & ( \Add1~89_sumout\ & ( (!\Selector10~4_combout\) # (((\R.aluOp.ALUOpSub~q\ & \Add2~89_sumout\)) # (\Selector10~1_combout\)) ) ) ) # ( \R.aluOp.ALUOpAdd~q\ 
-- & ( !\Add1~89_sumout\ & ( (!\Selector10~4_combout\) # (((\R.aluOp.ALUOpSub~q\ & \Add2~89_sumout\)) # (\Selector10~1_combout\)) ) ) ) # ( !\R.aluOp.ALUOpAdd~q\ & ( !\Add1~89_sumout\ & ( (!\Selector10~4_combout\) # (((\R.aluOp.ALUOpSub~q\ & 
-- \Add2~89_sumout\)) # (\Selector10~1_combout\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1011101110111111101110111011111110111011101111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector10~4_combout\,
	datab => \ALT_INV_Selector10~1_combout\,
	datac => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datad => \ALT_INV_Add2~89_sumout\,
	datae => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	dataf => \ALT_INV_Add1~89_sumout\,
	combout => \Selector10~5_combout\);

-- Location: FF_X77_Y2_N50
\R.aluRes[22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector10~5_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(22));

-- Location: LABCELL_X77_Y2_N3
\vAluRes~34\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~34_combout\ = ( \R.aluCalc~q\ & ( \Selector10~4_combout\ & ( !\Selector10~1_combout\ ) ) ) # ( !\R.aluCalc~q\ & ( \Selector10~4_combout\ & ( !\R.aluRes\(22) ) ) ) # ( !\R.aluCalc~q\ & ( !\Selector10~4_combout\ & ( !\R.aluRes\(22) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010101010101010000000000000000010101010101010101100110011001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluRes\(22),
	datab => \ALT_INV_Selector10~1_combout\,
	datae => \ALT_INV_R.aluCalc~q\,
	dataf => \ALT_INV_Selector10~4_combout\,
	combout => \vAluRes~34_combout\);

-- Location: MLABCELL_X78_Y2_N18
\vAluRes~19\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~19_combout\ = ( \Add1~89_sumout\ & ( \Add2~89_sumout\ & ( (!\vAluRes~34_combout\) # ((\R.aluCalc~q\ & ((\R.aluOp.ALUOpSub~q\) # (\R.aluOp.ALUOpAdd~q\)))) ) ) ) # ( !\Add1~89_sumout\ & ( \Add2~89_sumout\ & ( (!\vAluRes~34_combout\) # 
-- ((\R.aluOp.ALUOpSub~q\ & \R.aluCalc~q\)) ) ) ) # ( \Add1~89_sumout\ & ( !\Add2~89_sumout\ & ( (!\vAluRes~34_combout\) # ((\R.aluOp.ALUOpAdd~q\ & \R.aluCalc~q\)) ) ) ) # ( !\Add1~89_sumout\ & ( !\Add2~89_sumout\ & ( !\vAluRes~34_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111100000000111111110000010111111111000000111111111100000111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_R.aluCalc~q\,
	datad => \ALT_INV_vAluRes~34_combout\,
	datae => \ALT_INV_Add1~89_sumout\,
	dataf => \ALT_INV_Add2~89_sumout\,
	combout => \vAluRes~19_combout\);

-- Location: FF_X78_Y2_N19
\R.statusReg[0]_OTERM9_NEW_REG464\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \vAluRes~19_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.statusReg[0]_OTERM9_OTERM465\);

-- Location: LABCELL_X79_Y4_N18
\Equal3~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \Equal3~6_combout\ = ( \R.statusReg[0]_OTERM9_OTERM469\ & ( !\R.statusReg[0]_OTERM9_OTERM465\ & ( (\R.statusReg[0]_OTERM9_OTERM473\ & (!\R.statusReg[0]_OTERM9_OTERM467\ & (\R.statusReg[0]_OTERM9_OTERM471\ & !\R.statusReg[0]_OTERM9_OTERM463\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000001000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.statusReg[0]_OTERM9_OTERM473\,
	datab => \ALT_INV_R.statusReg[0]_OTERM9_OTERM467\,
	datac => \ALT_INV_R.statusReg[0]_OTERM9_OTERM471\,
	datad => \ALT_INV_R.statusReg[0]_OTERM9_OTERM463\,
	datae => \ALT_INV_R.statusReg[0]_OTERM9_OTERM469\,
	dataf => \ALT_INV_R.statusReg[0]_OTERM9_OTERM465\,
	combout => \Equal3~6_combout\);

-- Location: LABCELL_X74_Y6_N54
\ShiftLeft0~32\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~32_combout\ = ( \Mux234~0_combout\ & ( \Mux237~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((!\NxR.aluData2[0]~16_combout\)) # (\Mux235~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (((\Mux236~0_combout\) # 
-- (\NxR.aluData2[0]~16_combout\)))) ) ) ) # ( !\Mux234~0_combout\ & ( \Mux237~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (\Mux235~0_combout\ & (\NxR.aluData2[0]~16_combout\))) # (\NxR.aluData2[1]~17_combout\ & (((\Mux236~0_combout\) # 
-- (\NxR.aluData2[0]~16_combout\)))) ) ) ) # ( \Mux234~0_combout\ & ( !\Mux237~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((!\NxR.aluData2[0]~16_combout\)) # (\Mux235~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (((!\NxR.aluData2[0]~16_combout\ & 
-- \Mux236~0_combout\)))) ) ) ) # ( !\Mux234~0_combout\ & ( !\Mux237~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (\Mux235~0_combout\ & (\NxR.aluData2[0]~16_combout\))) # (\NxR.aluData2[1]~17_combout\ & (((!\NxR.aluData2[0]~16_combout\ & 
-- \Mux236~0_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001001010010101000101111001000000111010101111010011111110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datab => \ALT_INV_Mux235~0_combout\,
	datac => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datad => \ALT_INV_Mux236~0_combout\,
	datae => \ALT_INV_Mux234~0_combout\,
	dataf => \ALT_INV_Mux237~0_combout\,
	combout => \ShiftLeft0~32_combout\);

-- Location: FF_X74_Y6_N56
\ShiftLeft0~32_NEW_REG296\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~32_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~32_OTERM297\);

-- Location: LABCELL_X74_Y5_N12
\ShiftLeft0~40\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~40_combout\ = ( \NxR.aluData2[1]~17_combout\ & ( \Mux232~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\) # (\Mux233~0_combout\) ) ) ) # ( !\NxR.aluData2[1]~17_combout\ & ( \Mux232~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & 
-- (\Mux230~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & ((\Mux231~0_combout\))) ) ) ) # ( \NxR.aluData2[1]~17_combout\ & ( !\Mux232~0_combout\ & ( (\Mux233~0_combout\ & \NxR.aluData2[0]~16_combout\) ) ) ) # ( !\NxR.aluData2[1]~17_combout\ & ( 
-- !\Mux232~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (\Mux230~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & ((\Mux231~0_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000110000111111000100010001000100001100001111111101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux233~0_combout\,
	datab => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datac => \ALT_INV_Mux230~0_combout\,
	datad => \ALT_INV_Mux231~0_combout\,
	datae => \ALT_INV_NxR.aluData2[1]~17_combout\,
	dataf => \ALT_INV_Mux232~0_combout\,
	combout => \ShiftLeft0~40_combout\);

-- Location: FF_X74_Y5_N13
\ShiftLeft0~40_NEW_REG754\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~40_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~40_OTERM755\);

-- Location: LABCELL_X74_Y3_N30
\ShiftLeft0~49\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~49_combout\ = ( \NxR.aluData2[0]~16_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( \Mux229~0_combout\ ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( \Mux228~0_combout\ ) ) ) # ( \NxR.aluData2[0]~16_combout\ & ( 
-- !\NxR.aluData2[1]~17_combout\ & ( \Mux227~0_combout\ ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( !\NxR.aluData2[1]~17_combout\ & ( \Mux226~0_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111001100110011001100000000111111110101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux229~0_combout\,
	datab => \ALT_INV_Mux227~0_combout\,
	datac => \ALT_INV_Mux226~0_combout\,
	datad => \ALT_INV_Mux228~0_combout\,
	datae => \ALT_INV_NxR.aluData2[0]~16_combout\,
	dataf => \ALT_INV_NxR.aluData2[1]~17_combout\,
	combout => \ShiftLeft0~49_combout\);

-- Location: FF_X74_Y3_N31
\ShiftLeft0~49_NEW_REG760\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~49_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~49_OTERM761\);

-- Location: MLABCELL_X72_Y8_N54
\ShiftLeft0~50\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~50_combout\ = ( \ShiftLeft0~40_OTERM755\ & ( \ShiftLeft0~49_OTERM761\ & ( (!\R.aluData2\(3)) # ((!\R.aluData2\(2) & ((\ShiftLeft0~32_OTERM297\))) # (\R.aluData2\(2) & (\ShiftLeft0~24_OTERM293\))) ) ) ) # ( !\ShiftLeft0~40_OTERM755\ & ( 
-- \ShiftLeft0~49_OTERM761\ & ( (!\R.aluData2\(2) & (((!\R.aluData2\(3)) # (\ShiftLeft0~32_OTERM297\)))) # (\R.aluData2\(2) & (\ShiftLeft0~24_OTERM293\ & ((\R.aluData2\(3))))) ) ) ) # ( \ShiftLeft0~40_OTERM755\ & ( !\ShiftLeft0~49_OTERM761\ & ( 
-- (!\R.aluData2\(2) & (((\ShiftLeft0~32_OTERM297\ & \R.aluData2\(3))))) # (\R.aluData2\(2) & (((!\R.aluData2\(3))) # (\ShiftLeft0~24_OTERM293\))) ) ) ) # ( !\ShiftLeft0~40_OTERM755\ & ( !\ShiftLeft0~49_OTERM761\ & ( (\R.aluData2\(3) & ((!\R.aluData2\(2) & 
-- ((\ShiftLeft0~32_OTERM297\))) # (\R.aluData2\(2) & (\ShiftLeft0~24_OTERM293\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110101000011110011010111110000001101011111111100110101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~24_OTERM293\,
	datab => \ALT_INV_ShiftLeft0~32_OTERM297\,
	datac => \ALT_INV_R.aluData2\(2),
	datad => \ALT_INV_R.aluData2\(3),
	datae => \ALT_INV_ShiftLeft0~40_OTERM755\,
	dataf => \ALT_INV_ShiftLeft0~49_OTERM761\,
	combout => \ShiftLeft0~50_combout\);

-- Location: MLABCELL_X82_Y4_N18
\Selector4~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector4~0_combout\ = ( \R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( \R.aluOp.ALUOpOr~q\ & ( (!\R.aluData1\(28) & (!\R.aluData2\(28) & !\Selector17~0_OTERM391\)) ) ) ) # ( !\R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( \R.aluOp.ALUOpOr~q\ & ( (!\R.aluData1\(28) & 
-- (!\R.aluData2\(28) & !\Selector17~0_OTERM391\)) ) ) ) # ( \R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( !\R.aluOp.ALUOpOr~q\ & ( (!\Selector17~0_OTERM391\ & ((!\R.aluData1\(28) & ((!\R.aluData2\(28)) # (!\R.aluOp.ALUOpXor~DUPLICATE_q\))) # (\R.aluData1\(28) & 
-- (!\R.aluData2\(28) & !\R.aluOp.ALUOpXor~DUPLICATE_q\)))) ) ) ) # ( !\R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( !\R.aluOp.ALUOpOr~q\ & ( (!\Selector17~0_OTERM391\ & ((!\R.aluOp.ALUOpXor~DUPLICATE_q\) # (!\R.aluData1\(28) $ (\R.aluData2\(28))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111000010010000111000001000000010000000100000001000000010000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData1\(28),
	datab => \ALT_INV_R.aluData2\(28),
	datac => \ALT_INV_Selector17~0_OTERM391\,
	datad => \ALT_INV_R.aluOp.ALUOpXor~DUPLICATE_q\,
	datae => \ALT_INV_R.aluOp.ALUOpAnd~DUPLICATE_q\,
	dataf => \ALT_INV_R.aluOp.ALUOpOr~q\,
	combout => \Selector4~0_combout\);

-- Location: MLABCELL_X78_Y4_N36
\Selector20~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector20~5_combout\ = ( \ShiftRight1~3_OTERM13\ & ( (!\Selector20~0_OTERM769\ & ((!\Selector31~0_OTERM349\) # (\ShiftRight0~7_OTERM233DUPLICATE_q\))) ) ) # ( !\ShiftRight1~3_OTERM13\ & ( !\Selector20~0_OTERM769\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111100000000111111110000000011001111000000001100111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Selector31~0_OTERM349\,
	datac => \ALT_INV_ShiftRight0~7_OTERM233DUPLICATE_q\,
	datad => \ALT_INV_Selector20~0_OTERM769\,
	dataf => \ALT_INV_ShiftRight1~3_OTERM13\,
	combout => \Selector20~5_combout\);

-- Location: MLABCELL_X78_Y4_N42
\Selector4~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector4~1_combout\ = ( \Selector20~5_combout\ & ( \R.aluOp.ALUOpSLL~q\ & ( (!\Selector4~0_combout\) # ((!\R.aluData2\(4) & ((\ShiftLeft0~50_combout\))) # (\R.aluData2\(4) & (\ShiftLeft0~17_combout\))) ) ) ) # ( !\Selector20~5_combout\ & ( 
-- \R.aluOp.ALUOpSLL~q\ & ( (!\R.aluData2\(4)) # ((!\Selector4~0_combout\) # (\ShiftLeft0~17_combout\)) ) ) ) # ( \Selector20~5_combout\ & ( !\R.aluOp.ALUOpSLL~q\ & ( !\Selector4~0_combout\ ) ) ) # ( !\Selector20~5_combout\ & ( !\R.aluOp.ALUOpSLL~q\ & ( 
-- (!\R.aluData2\(4)) # (!\Selector4~0_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111110101010111111110000000011111111101110111111111100011011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(4),
	datab => \ALT_INV_ShiftLeft0~17_combout\,
	datac => \ALT_INV_ShiftLeft0~50_combout\,
	datad => \ALT_INV_Selector4~0_combout\,
	datae => \ALT_INV_Selector20~5_combout\,
	dataf => \ALT_INV_R.aluOp.ALUOpSLL~q\,
	combout => \Selector4~1_combout\);

-- Location: LABCELL_X79_Y5_N24
\Add2~113\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~113_sumout\ = SUM(( !\R.aluData1\(28) $ (\R.aluData2\(28)) ) + ( \Add2~111\ ) + ( \Add2~110\ ))
-- \Add2~114\ = CARRY(( !\R.aluData1\(28) $ (\R.aluData2\(28)) ) + ( \Add2~111\ ) + ( \Add2~110\ ))
-- \Add2~115\ = SHARE((\R.aluData1\(28) & !\R.aluData2\(28)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000001100110000000000000000000000001100110000110011",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluData1\(28),
	datad => \ALT_INV_R.aluData2\(28),
	cin => \Add2~110\,
	sharein => \Add2~111\,
	sumout => \Add2~113_sumout\,
	cout => \Add2~114\,
	shareout => \Add2~115\);

-- Location: MLABCELL_X78_Y4_N51
\Selector4~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector4~2_combout\ = ( \Add2~113_sumout\ & ( (((\R.aluOp.ALUOpAdd~q\ & \Add1~113_sumout\)) # (\R.aluOp.ALUOpSub~q\)) # (\Selector4~1_combout\) ) ) # ( !\Add2~113_sumout\ & ( ((\R.aluOp.ALUOpAdd~q\ & \Add1~113_sumout\)) # (\Selector4~1_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001111100011111000111110001111100011111111111110001111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datab => \ALT_INV_Add1~113_sumout\,
	datac => \ALT_INV_Selector4~1_combout\,
	datad => \ALT_INV_R.aluOp.ALUOpSub~q\,
	dataf => \ALT_INV_Add2~113_sumout\,
	combout => \Selector4~2_combout\);

-- Location: FF_X78_Y4_N53
\R.aluRes[28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector4~2_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(28));

-- Location: MLABCELL_X78_Y4_N54
\vAluRes~48\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~48_combout\ = ( !\R.aluCalc~q\ & ( (((\R.aluRes\(28)))) ) ) # ( \R.aluCalc~q\ & ( ((!\R.aluOp.ALUOpSub~q\ & (\R.aluOp.ALUOpAdd~q\ & (\Add1~113_sumout\))) # (\R.aluOp.ALUOpSub~q\ & (((\R.aluOp.ALUOpAdd~q\ & \Add1~113_sumout\)) # 
-- (\Add2~113_sumout\)))) # (\Selector4~1_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100001111001100110011111100001111000011110111011101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datab => \ALT_INV_Selector4~1_combout\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_Add1~113_sumout\,
	datae => \ALT_INV_R.aluCalc~q\,
	dataf => \ALT_INV_Add2~113_sumout\,
	datag => \ALT_INV_R.aluRes\(28),
	combout => \vAluRes~48_combout\);

-- Location: FF_X78_Y4_N56
\R.statusReg[0]_NEW_REG4\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \vAluRes~48_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.statusReg[0]_OTERM5\);

-- Location: FF_X79_Y5_N34
\R.statusReg[0]_OTERM7_NEW_REG490\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Add2~125_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.statusReg[0]_OTERM7_OTERM491\);

-- Location: LABCELL_X77_Y8_N48
\ShiftLeft0~23\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~23_combout\ = ( \ShiftLeft0~9_OTERM461\ & ( \R.aluData2\(3) & ( (!\R.aluData2\(2)) # (\ShiftLeft0~3_OTERM223\) ) ) ) # ( !\ShiftLeft0~9_OTERM461\ & ( \R.aluData2\(3) & ( (\R.aluData2\(2) & \ShiftLeft0~3_OTERM223\) ) ) ) # ( 
-- \ShiftLeft0~9_OTERM461\ & ( !\R.aluData2\(3) & ( (!\R.aluData2\(2) & ((\ShiftLeft0~22_OTERM737\))) # (\R.aluData2\(2) & (\ShiftLeft0~14_OTERM753\)) ) ) ) # ( !\ShiftLeft0~9_OTERM461\ & ( !\R.aluData2\(3) & ( (!\R.aluData2\(2) & 
-- ((\ShiftLeft0~22_OTERM737\))) # (\R.aluData2\(2) & (\ShiftLeft0~14_OTERM753\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001110100011101000111010001110100000000001100111100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~14_OTERM753\,
	datab => \ALT_INV_R.aluData2\(2),
	datac => \ALT_INV_ShiftLeft0~22_OTERM737\,
	datad => \ALT_INV_ShiftLeft0~3_OTERM223\,
	datae => \ALT_INV_ShiftLeft0~9_OTERM461\,
	dataf => \ALT_INV_R.aluData2\(3),
	combout => \ShiftLeft0~23_combout\);

-- Location: MLABCELL_X72_Y5_N39
\Selector1~0_RTM0773\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector1~0_RTM0773_combout\ = ( \NxR.aluData2[31]~29_combout\ & ( \R.aluOp.ALUOpSRA_OTERM363\ & ( ((\Mux223~0_combout\) # (\R.aluOp.ALUOpXor_OTERM355\)) # (\R.aluOp.ALUOpOr_OTERM353\) ) ) ) # ( !\NxR.aluData2[31]~29_combout\ & ( 
-- \R.aluOp.ALUOpSRA_OTERM363\ & ( \Mux223~0_combout\ ) ) ) # ( \NxR.aluData2[31]~29_combout\ & ( !\R.aluOp.ALUOpSRA_OTERM363\ & ( ((!\Mux223~0_combout\ & (\R.aluOp.ALUOpXor_OTERM355\)) # (\Mux223~0_combout\ & ((\R.aluOp.ALUOpAnd_OTERM357\)))) # 
-- (\R.aluOp.ALUOpOr_OTERM353\) ) ) ) # ( !\NxR.aluData2[31]~29_combout\ & ( !\R.aluOp.ALUOpSRA_OTERM363\ & ( (\Mux223~0_combout\ & ((\R.aluOp.ALUOpXor_OTERM355\) # (\R.aluOp.ALUOpOr_OTERM353\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001110111011101110101111100000000111111110111011111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpOr_OTERM353\,
	datab => \ALT_INV_R.aluOp.ALUOpXor_OTERM355\,
	datac => \ALT_INV_R.aluOp.ALUOpAnd_OTERM357\,
	datad => \ALT_INV_Mux223~0_combout\,
	datae => \ALT_INV_NxR.aluData2[31]~29_combout\,
	dataf => \ALT_INV_R.aluOp.ALUOpSRA_OTERM363\,
	combout => \Selector1~0_RTM0773_combout\);

-- Location: FF_X72_Y5_N40
\Selector1~0_NEW_REG770\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector1~0_RTM0773_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector1~0_OTERM771\);

-- Location: LABCELL_X77_Y7_N21
\Selector1~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector1~1_combout\ = ( \R.aluData2\(4) & ( !\Selector1~0_OTERM771\ ) ) # ( !\R.aluData2\(4) & ( (!\Selector1~0_OTERM771\ & ((!\ShiftRight0~4_OTERM31\) # ((!\R.aluOp.ALUOpSRL~q\) # (\ShiftRight0~7_OTERM233DUPLICATE_q\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111101100000000111110110000000011111111000000001111111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight0~4_OTERM31\,
	datab => \ALT_INV_ShiftRight0~7_OTERM233DUPLICATE_q\,
	datac => \ALT_INV_R.aluOp.ALUOpSRL~q\,
	datad => \ALT_INV_Selector1~0_OTERM771\,
	dataf => \ALT_INV_R.aluData2\(4),
	combout => \Selector1~1_combout\);

-- Location: LABCELL_X73_Y5_N24
\ShiftLeft0~55\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~55_combout\ = ( \NxR.aluData2[0]~16_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( \Mux226~0_combout\ ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( \Mux225~0_combout\ ) ) ) # ( \NxR.aluData2[0]~16_combout\ & ( 
-- !\NxR.aluData2[1]~17_combout\ & ( \Mux224~0_combout\ ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( !\NxR.aluData2[1]~17_combout\ & ( \Mux223~0_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110011000000001111111101010101010101010000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux225~0_combout\,
	datab => \ALT_INV_Mux223~0_combout\,
	datac => \ALT_INV_Mux226~0_combout\,
	datad => \ALT_INV_Mux224~0_combout\,
	datae => \ALT_INV_NxR.aluData2[0]~16_combout\,
	dataf => \ALT_INV_NxR.aluData2[1]~17_combout\,
	combout => \ShiftLeft0~55_combout\);

-- Location: FF_X73_Y5_N25
\ShiftLeft0~55_NEW_REG766\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~55_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~55_OTERM767\);

-- Location: LABCELL_X79_Y7_N18
\ShiftLeft0~56\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~56_combout\ = ( \ShiftLeft0~38_OTERM789\ & ( \R.aluData2\(3) & ( (!\R.aluData2\(2)) # (\ShiftLeft0~30_OTERM601\) ) ) ) # ( !\ShiftLeft0~38_OTERM789\ & ( \R.aluData2\(3) & ( (\R.aluData2\(2) & \ShiftLeft0~30_OTERM601\) ) ) ) # ( 
-- \ShiftLeft0~38_OTERM789\ & ( !\R.aluData2\(3) & ( (!\R.aluData2\(2) & ((\ShiftLeft0~55_OTERM767\))) # (\R.aluData2\(2) & (\ShiftLeft0~47_OTERM759\)) ) ) ) # ( !\ShiftLeft0~38_OTERM789\ & ( !\R.aluData2\(3) & ( (!\R.aluData2\(2) & 
-- ((\ShiftLeft0~55_OTERM767\))) # (\R.aluData2\(2) & (\ShiftLeft0~47_OTERM759\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000110111011000100011011101100000101000001011010111110101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(2),
	datab => \ALT_INV_ShiftLeft0~47_OTERM759\,
	datac => \ALT_INV_ShiftLeft0~30_OTERM601\,
	datad => \ALT_INV_ShiftLeft0~55_OTERM767\,
	datae => \ALT_INV_ShiftLeft0~38_OTERM789\,
	dataf => \ALT_INV_R.aluData2\(3),
	combout => \ShiftLeft0~56_combout\);

-- Location: LABCELL_X79_Y7_N36
\Selector1~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector1~2_combout\ = ( \Selector1~1_combout\ & ( \ShiftLeft0~56_combout\ & ( (\R.aluOp.ALUOpSLL~q\ & ((!\R.aluData2\(4)) # (\ShiftLeft0~23_combout\))) ) ) ) # ( !\Selector1~1_combout\ & ( \ShiftLeft0~56_combout\ ) ) # ( \Selector1~1_combout\ & ( 
-- !\ShiftLeft0~56_combout\ & ( (\R.aluData2\(4) & (\ShiftLeft0~23_combout\ & \R.aluOp.ALUOpSLL~q\)) ) ) ) # ( !\Selector1~1_combout\ & ( !\ShiftLeft0~56_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111000000000000010111111111111111110000000010101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(4),
	datac => \ALT_INV_ShiftLeft0~23_combout\,
	datad => \ALT_INV_R.aluOp.ALUOpSLL~q\,
	datae => \ALT_INV_Selector1~1_combout\,
	dataf => \ALT_INV_ShiftLeft0~56_combout\,
	combout => \Selector1~2_combout\);

-- Location: FF_X79_Y7_N4
\R.statusReg[0]_OTERM7_NEW_REG480\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Selector1~2_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.statusReg[0]_OTERM7_OTERM481\);

-- Location: FF_X79_Y5_N52
\R.statusReg[0]_OTERM7_NEW_REG482\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \vAluRes~25_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.statusReg[0]_OTERM7_OTERM483\);

-- Location: LABCELL_X83_Y7_N24
\Equal3~19\ : cyclonev_lcell_comb
-- Equation(s):
-- \Equal3~19_combout\ = ( \Selector1~2_combout\ & ( \R.aluCalc~q\ ) ) # ( !\Selector1~2_combout\ & ( (\R.aluCalc~q\ & \R.aluOp.ALUOpSub~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101010101010101010100000101000001010101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datae => \ALT_INV_Selector1~2_combout\,
	combout => \Equal3~19_combout\);

-- Location: FF_X83_Y7_N25
\R.statusReg[0]_OTERM7_NEW_REG488\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Equal3~19_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.statusReg[0]_OTERM7_OTERM489\);

-- Location: MLABCELL_X78_Y5_N33
\Add1~125\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~125_sumout\ = SUM(( \R.aluData2\(31) ) + ( \R.aluData1\(31) ) + ( \Add1~122\ ))
-- \Add1~126\ = CARRY(( \R.aluData2\(31) ) + ( \R.aluData1\(31) ) + ( \Add1~122\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluData2\(31),
	datac => \ALT_INV_R.aluData1\(31),
	cin => \Add1~122\,
	sumout => \Add1~125_sumout\,
	cout => \Add1~126\);

-- Location: MLABCELL_X78_Y5_N9
\Add1~93\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~93_sumout\ = SUM(( \R.aluData2\(23) ) + ( \R.aluData1\(23) ) + ( \Add1~90\ ))
-- \Add1~94\ = CARRY(( \R.aluData2\(23) ) + ( \R.aluData1\(23) ) + ( \Add1~90\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluData1\(23),
	datad => \ALT_INV_R.aluData2\(23),
	cin => \Add1~90\,
	sumout => \Add1~93_sumout\,
	cout => \Add1~94\);

-- Location: MLABCELL_X78_Y5_N12
\Add1~97\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~97_sumout\ = SUM(( \R.aluData2\(24) ) + ( \R.aluData1\(24) ) + ( \Add1~94\ ))
-- \Add1~98\ = CARRY(( \R.aluData2\(24) ) + ( \R.aluData1\(24) ) + ( \Add1~94\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluData1\(24),
	datad => \ALT_INV_R.aluData2\(24),
	cin => \Add1~94\,
	sumout => \Add1~97_sumout\,
	cout => \Add1~98\);

-- Location: MLABCELL_X78_Y5_N15
\Add1~101\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~101_sumout\ = SUM(( \R.aluData2[25]~DUPLICATE_q\ ) + ( \R.aluData1\(25) ) + ( \Add1~98\ ))
-- \Add1~102\ = CARRY(( \R.aluData2[25]~DUPLICATE_q\ ) + ( \R.aluData1\(25) ) + ( \Add1~98\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData1\(25),
	datab => \ALT_INV_R.aluData2[25]~DUPLICATE_q\,
	cin => \Add1~98\,
	sumout => \Add1~101_sumout\,
	cout => \Add1~102\);

-- Location: MLABCELL_X82_Y5_N0
\Selector7~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector7~3_combout\ = ( \Selector7~5_combout\ & ( \R.aluOp.ALUOpSub~q\ ) ) # ( !\Selector7~5_combout\ & ( \R.aluOp.ALUOpSub~q\ & ( (((\R.aluOp.ALUOpAdd~q\ & \Add1~101_sumout\)) # (\Selector7~1_combout\)) # (\Add2~101_sumout\) ) ) ) # ( 
-- \Selector7~5_combout\ & ( !\R.aluOp.ALUOpSub~q\ ) ) # ( !\Selector7~5_combout\ & ( !\R.aluOp.ALUOpSub~q\ & ( ((\R.aluOp.ALUOpAdd~q\ & \Add1~101_sumout\)) # (\Selector7~1_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111101011111111111111111111100111111011111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datab => \ALT_INV_Add2~101_sumout\,
	datac => \ALT_INV_Selector7~1_combout\,
	datad => \ALT_INV_Add1~101_sumout\,
	datae => \ALT_INV_Selector7~5_combout\,
	dataf => \ALT_INV_R.aluOp.ALUOpSub~q\,
	combout => \Selector7~3_combout\);

-- Location: FF_X82_Y5_N2
\R.aluRes[25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector7~3_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(25));

-- Location: LABCELL_X83_Y3_N30
\vAluRes~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~26_combout\ = ( \R.aluRes\(25) & ( !\R.aluCalc~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datae => \ALT_INV_R.aluRes\(25),
	dataf => \ALT_INV_R.aluCalc~q\,
	combout => \vAluRes~26_combout\);

-- Location: LABCELL_X77_Y3_N12
\Equal3~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Equal3~18_combout\ = ( \Add1~125_sumout\ & ( !\vAluRes~26_combout\ & ( (!\vAluRes~30_combout\ & (!\vAluRes~28_combout\ & ((!\R.aluOp.ALUOpAdd~q\) # (!\R.aluCalc~q\)))) ) ) ) # ( !\Add1~125_sumout\ & ( !\vAluRes~26_combout\ & ( (!\vAluRes~30_combout\ & 
-- !\vAluRes~28_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1100110000000000110010000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datab => \ALT_INV_vAluRes~30_combout\,
	datac => \ALT_INV_R.aluCalc~q\,
	datad => \ALT_INV_vAluRes~28_combout\,
	datae => \ALT_INV_Add1~125_sumout\,
	dataf => \ALT_INV_vAluRes~26_combout\,
	combout => \Equal3~18_combout\);

-- Location: FF_X77_Y3_N13
\R.statusReg[0]_OTERM7_NEW_REG486\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Equal3~18_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.statusReg[0]_OTERM7_OTERM487\);

-- Location: MLABCELL_X78_Y5_N18
\Add1~105\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~105_sumout\ = SUM(( \R.aluData1\(26) ) + ( \R.aluData2\(26) ) + ( \Add1~102\ ))
-- \Add1~106\ = CARRY(( \R.aluData1\(26) ) + ( \R.aluData2\(26) ) + ( \Add1~102\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluData2\(26),
	datad => \ALT_INV_R.aluData1\(26),
	cin => \Add1~102\,
	sumout => \Add1~105_sumout\,
	cout => \Add1~106\);

-- Location: MLABCELL_X78_Y7_N36
\vAluRes~27\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~27_combout\ = ( \Add2~105_sumout\ & ( \R.aluCalc~q\ & ( (!\Selector6~1_combout\) # (((\R.aluOp.ALUOpAdd~q\ & \Add1~105_sumout\)) # (\R.aluOp.ALUOpSub~q\)) ) ) ) # ( !\Add2~105_sumout\ & ( \R.aluCalc~q\ & ( (!\Selector6~1_combout\) # 
-- ((\R.aluOp.ALUOpAdd~q\ & \Add1~105_sumout\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000010101010101110111010111110111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector6~1_combout\,
	datab => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datac => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datad => \ALT_INV_Add1~105_sumout\,
	datae => \ALT_INV_Add2~105_sumout\,
	dataf => \ALT_INV_R.aluCalc~q\,
	combout => \vAluRes~27_combout\);

-- Location: FF_X78_Y7_N37
\R.statusReg[0]_OTERM7_NEW_REG484\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \vAluRes~27_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.statusReg[0]_OTERM7_OTERM485\);

-- Location: LABCELL_X80_Y7_N54
\Equal3~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Equal3~2_combout\ = ( \R.statusReg[0]_OTERM7_OTERM487\ & ( !\R.statusReg[0]_OTERM7_OTERM485\ & ( (!\R.statusReg[0]_OTERM7_OTERM483\ & ((!\R.statusReg[0]_OTERM7_OTERM489\) # ((!\R.statusReg[0]_OTERM7_OTERM491\ & !\R.statusReg[0]_OTERM7_OTERM481\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.statusReg[0]_OTERM7_OTERM491\,
	datab => \ALT_INV_R.statusReg[0]_OTERM7_OTERM481\,
	datac => \ALT_INV_R.statusReg[0]_OTERM7_OTERM483\,
	datad => \ALT_INV_R.statusReg[0]_OTERM7_OTERM489\,
	datae => \ALT_INV_R.statusReg[0]_OTERM7_OTERM487\,
	dataf => \ALT_INV_R.statusReg[0]_OTERM7_OTERM485\,
	combout => \Equal3~2_combout\);

-- Location: MLABCELL_X78_Y8_N3
\vAluRes~33\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~33_combout\ = (!\R.aluCalc~q\ & (!\R.aluRes\(20))) # (\R.aluCalc~q\ & (((\Selector12~4_combout\ & !\Selector12~1_combout\))))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000101110001000100010111000100010001011100010001000101110001000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluRes\(20),
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_Selector12~4_combout\,
	datad => \ALT_INV_Selector12~1_combout\,
	combout => \vAluRes~33_combout\);

-- Location: LABCELL_X79_Y8_N42
\vAluRes~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~17_combout\ = ( \R.aluCalc~q\ & ( \Add1~81_sumout\ & ( ((!\vAluRes~33_combout\) # ((\Add2~81_sumout\ & \R.aluOp.ALUOpSub~q\))) # (\R.aluOp.ALUOpAdd~q\) ) ) ) # ( !\R.aluCalc~q\ & ( \Add1~81_sumout\ & ( !\vAluRes~33_combout\ ) ) ) # ( 
-- \R.aluCalc~q\ & ( !\Add1~81_sumout\ & ( (!\vAluRes~33_combout\) # ((\Add2~81_sumout\ & \R.aluOp.ALUOpSub~q\)) ) ) ) # ( !\R.aluCalc~q\ & ( !\Add1~81_sumout\ & ( !\vAluRes~33_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111100000000111111110000001111111111000000001111111101010111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datab => \ALT_INV_Add2~81_sumout\,
	datac => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datad => \ALT_INV_vAluRes~33_combout\,
	datae => \ALT_INV_R.aluCalc~q\,
	dataf => \ALT_INV_Add1~81_sumout\,
	combout => \vAluRes~17_combout\);

-- Location: FF_X80_Y5_N22
\R.aluRes[0]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector32~8_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes[0]~DUPLICATE_q\);

-- Location: LABCELL_X80_Y5_N30
\vAluRes~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~0_combout\ = ( \R.aluCalc~q\ & ( \Selector32~1_combout\ ) ) # ( !\R.aluCalc~q\ & ( \Selector32~1_combout\ & ( \R.aluRes[0]~DUPLICATE_q\ ) ) ) # ( \R.aluCalc~q\ & ( !\Selector32~1_combout\ & ( !\Selector32~7_combout\ ) ) ) # ( !\R.aluCalc~q\ & ( 
-- !\Selector32~1_combout\ & ( \R.aluRes[0]~DUPLICATE_q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110011111100001111000000110011001100111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluRes[0]~DUPLICATE_q\,
	datac => \ALT_INV_Selector32~7_combout\,
	datae => \ALT_INV_R.aluCalc~q\,
	dataf => \ALT_INV_Selector32~1_combout\,
	combout => \vAluRes~0_combout\);

-- Location: LABCELL_X79_Y8_N6
\Equal3~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Equal3~1_combout\ = ( !\vAluRes~8_combout\ & ( !\vAluRes~0_combout\ & ( (!\vAluRes~1_combout\ & (!\vAluRes~17_combout\ & (!\vAluRes~56_combout\ & !\vAluRes~2_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000000000000000000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluRes~1_combout\,
	datab => \ALT_INV_vAluRes~17_combout\,
	datac => \ALT_INV_vAluRes~56_combout\,
	datad => \ALT_INV_vAluRes~2_combout\,
	datae => \ALT_INV_vAluRes~8_combout\,
	dataf => \ALT_INV_vAluRes~0_combout\,
	combout => \Equal3~1_combout\);

-- Location: FF_X79_Y8_N7
\R.statusReg[0]_OTERM11_NEW_REG374\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Equal3~1_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.statusReg[0]_OTERM11_OTERM375\);

-- Location: FF_X80_Y4_N7
\R.statusReg[0]_OTERM11_NEW_REG370\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector9~5_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.statusReg[0]_OTERM11_OTERM371\);

-- Location: FF_X79_Y3_N43
\R.statusReg[0]_OTERM11_NEW_REG368\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector14~3_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.statusReg[0]_OTERM11_OTERM369\);

-- Location: FF_X80_Y4_N37
\R.statusReg[0]_OTERM11_NEW_REG372\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector8~4_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.statusReg[0]_OTERM11_OTERM373\);

-- Location: FF_X84_Y4_N2
\R.statusReg[0]_OTERM11_NEW_REG366\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.aluCalc~q\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.statusReg[0]_OTERM11_OTERM367\);

-- Location: LABCELL_X73_Y8_N6
\Selector23~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector23~1_combout\ = ( \ShiftLeft0~1_OTERM255\ & ( \R.aluData2\(3) & ( (!\R.aluData2\(2) & \Selector27~0_OTERM385\) ) ) ) # ( \ShiftLeft0~1_OTERM255\ & ( !\R.aluData2\(3) & ( (\Selector27~0_OTERM385\ & ((!\R.aluData2\(2) & 
-- ((\ShiftLeft0~12_OTERM791\))) # (\R.aluData2\(2) & (\ShiftLeft0~7_OTERM205\)))) ) ) ) # ( !\ShiftLeft0~1_OTERM255\ & ( !\R.aluData2\(3) & ( (\Selector27~0_OTERM385\ & ((!\R.aluData2\(2) & ((\ShiftLeft0~12_OTERM791\))) # (\R.aluData2\(2) & 
-- (\ShiftLeft0~7_OTERM205\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110101000000000011010100000000000000000000000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~7_OTERM205\,
	datab => \ALT_INV_ShiftLeft0~12_OTERM791\,
	datac => \ALT_INV_R.aluData2\(2),
	datad => \ALT_INV_Selector27~0_OTERM385\,
	datae => \ALT_INV_ShiftLeft0~1_OTERM255\,
	dataf => \ALT_INV_R.aluData2\(3),
	combout => \Selector23~1_combout\);

-- Location: LABCELL_X77_Y9_N48
\Selector23~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector23~2_combout\ = ( \ShiftRight1~12_OTERM57\ & ( \ShiftRight1~13_OTERM15\ & ( (\Selector31~6_OTERM381\ & ((!\R.aluData2\(3)) # (\R.aluData1\(31)))) ) ) ) # ( !\ShiftRight1~12_OTERM57\ & ( \ShiftRight1~13_OTERM15\ & ( (\Selector31~6_OTERM381\ & 
-- ((!\R.aluData2\(3) & ((\R.aluData2\(2)))) # (\R.aluData2\(3) & (\R.aluData1\(31))))) ) ) ) # ( \ShiftRight1~12_OTERM57\ & ( !\ShiftRight1~13_OTERM15\ & ( (\Selector31~6_OTERM381\ & ((!\R.aluData2\(3) & ((!\R.aluData2\(2)))) # (\R.aluData2\(3) & 
-- (\R.aluData1\(31))))) ) ) ) # ( !\ShiftRight1~12_OTERM57\ & ( !\ShiftRight1~13_OTERM15\ & ( (\R.aluData1\(31) & (\R.aluData2\(3) & \Selector31~6_OTERM381\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000101000000001100010100000000001101010000000011110101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData1\(31),
	datab => \ALT_INV_R.aluData2\(2),
	datac => \ALT_INV_R.aluData2\(3),
	datad => \ALT_INV_Selector31~6_OTERM381\,
	datae => \ALT_INV_ShiftRight1~12_OTERM57\,
	dataf => \ALT_INV_ShiftRight1~13_OTERM15\,
	combout => \Selector23~2_combout\);

-- Location: LABCELL_X74_Y7_N39
\Selector23~3_RTM0425\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector23~3_RTM0425_combout\ = ( \R.aluOp.ALUOpAnd_OTERM357\ & ( (!\Mux245~0_combout\ & (\NxR.aluData2[9]~12_combout\ & ((\R.aluOp.ALUOpXor_OTERM355\) # (\R.aluOp.ALUOpOr_OTERM353\)))) # (\Mux245~0_combout\ & (((\NxR.aluData2[9]~12_combout\) # 
-- (\R.aluOp.ALUOpXor_OTERM355\)) # (\R.aluOp.ALUOpOr_OTERM353\))) ) ) # ( !\R.aluOp.ALUOpAnd_OTERM357\ & ( (!\R.aluOp.ALUOpOr_OTERM353\ & (\R.aluOp.ALUOpXor_OTERM355\ & (!\Mux245~0_combout\ $ (!\NxR.aluData2[9]~12_combout\)))) # (\R.aluOp.ALUOpOr_OTERM353\ 
-- & (((\NxR.aluData2[9]~12_combout\)) # (\Mux245~0_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001001101011101000100110101110100010011011111110001001101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpOr_OTERM353\,
	datab => \ALT_INV_Mux245~0_combout\,
	datac => \ALT_INV_R.aluOp.ALUOpXor_OTERM355\,
	datad => \ALT_INV_NxR.aluData2[9]~12_combout\,
	dataf => \ALT_INV_R.aluOp.ALUOpAnd_OTERM357\,
	combout => \Selector23~3_RTM0425_combout\);

-- Location: FF_X74_Y7_N40
\Selector23~3_NEW_REG422\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector23~3_RTM0425_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector23~3_OTERM423\);

-- Location: LABCELL_X77_Y9_N6
\Selector23~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector23~4_combout\ = ( \Selector31~7_OTERM383\ & ( \R.aluData2\(2) & ( (!\Selector23~3_OTERM423\ & ((!\ShiftRight0~0_OTERM17\) # (\R.aluData2\(3)))) ) ) ) # ( !\Selector31~7_OTERM383\ & ( \R.aluData2\(2) & ( !\Selector23~3_OTERM423\ ) ) ) # ( 
-- \Selector31~7_OTERM383\ & ( !\R.aluData2\(2) & ( (!\Selector23~3_OTERM423\ & ((!\ShiftRight1~12_OTERM57\) # (\R.aluData2\(3)))) ) ) ) # ( !\Selector31~7_OTERM383\ & ( !\R.aluData2\(2) & ( !\Selector23~3_OTERM423\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1100110011001100110011000100010011001100110011001100010011000100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(3),
	datab => \ALT_INV_Selector23~3_OTERM423\,
	datac => \ALT_INV_ShiftRight0~0_OTERM17\,
	datad => \ALT_INV_ShiftRight1~12_OTERM57\,
	datae => \ALT_INV_Selector31~7_OTERM383\,
	dataf => \ALT_INV_R.aluData2\(2),
	combout => \Selector23~4_combout\);

-- Location: LABCELL_X79_Y9_N18
\Selector23~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector23~7_combout\ = ( \Selector23~4_combout\ & ( \ShiftRight1~47_combout\ & ( (!\Selector23~2_combout\ & !\Selector31~5_OTERM599\) ) ) ) # ( \Selector23~4_combout\ & ( !\ShiftRight1~47_combout\ & ( !\Selector23~2_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000001010000010100000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector23~2_combout\,
	datac => \ALT_INV_Selector31~5_OTERM599\,
	datae => \ALT_INV_Selector23~4_combout\,
	dataf => \ALT_INV_ShiftRight1~47_combout\,
	combout => \Selector23~7_combout\);

-- Location: LABCELL_X80_Y3_N42
\Selector23~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector23~6_combout\ = ( \Add2~37_sumout\ & ( \Selector23~7_combout\ & ( (((\Add1~37_sumout\ & \R.aluOp.ALUOpAdd~q\)) # (\Selector23~1_combout\)) # (\R.aluOp.ALUOpSub~q\) ) ) ) # ( !\Add2~37_sumout\ & ( \Selector23~7_combout\ & ( ((\Add1~37_sumout\ & 
-- \R.aluOp.ALUOpAdd~q\)) # (\Selector23~1_combout\) ) ) ) # ( \Add2~37_sumout\ & ( !\Selector23~7_combout\ ) ) # ( !\Add2~37_sumout\ & ( !\Selector23~7_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111111111111111111100010001111111110001111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add1~37_sumout\,
	datab => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datac => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datad => \ALT_INV_Selector23~1_combout\,
	datae => \ALT_INV_Add2~37_sumout\,
	dataf => \ALT_INV_Selector23~7_combout\,
	combout => \Selector23~6_combout\);

-- Location: FF_X80_Y3_N44
\R.aluRes[9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector23~6_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(9));

-- Location: LABCELL_X80_Y3_N27
\Selector18~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector18~5_combout\ = ( \Selector18~3_combout\ & ( (!\R.aluOp.ALUOpSub~q\ & (\R.aluOp.ALUOpAdd~q\ & (\Add1~57_sumout\))) # (\R.aluOp.ALUOpSub~q\ & (((\R.aluOp.ALUOpAdd~q\ & \Add1~57_sumout\)) # (\Add2~57_sumout\))) ) ) # ( !\Selector18~3_combout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111111111111111111100000011010101110000001101010111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datab => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datac => \ALT_INV_Add1~57_sumout\,
	datad => \ALT_INV_Add2~57_sumout\,
	dataf => \ALT_INV_Selector18~3_combout\,
	combout => \Selector18~5_combout\);

-- Location: FF_X80_Y3_N28
\R.aluRes[14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector18~5_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(14));

-- Location: LABCELL_X80_Y3_N51
\Equal3~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \Equal3~11_combout\ = ( \R.aluRes\(14) & ( (\R.aluCalc~q\ & ((!\R.aluOp.ALUOpAdd~q\) # (!\Add1~57_sumout\))) ) ) # ( !\R.aluRes\(14) & ( (!\R.aluCalc~q\ & (!\R.aluRes\(9))) # (\R.aluCalc~q\ & (((!\R.aluOp.ALUOpAdd~q\) # (!\Add1~57_sumout\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1101110111011000110111011101100001010101010100000101010101010000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluCalc~q\,
	datab => \ALT_INV_R.aluRes\(9),
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_Add1~57_sumout\,
	dataf => \ALT_INV_R.aluRes\(14),
	combout => \Equal3~11_combout\);

-- Location: LABCELL_X80_Y3_N12
\Equal3~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \Equal3~7_combout\ = ( \Selector23~6_combout\ & ( \Equal3~11_combout\ & ( !\R.aluCalc~q\ ) ) ) # ( !\Selector23~6_combout\ & ( \Equal3~11_combout\ & ( (!\R.aluCalc~q\) # ((\Selector18~3_combout\ & ((!\R.aluOp.ALUOpSub~q\) # (!\Add2~57_sumout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011001100111111101100110011001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_Add2~57_sumout\,
	datad => \ALT_INV_Selector18~3_combout\,
	datae => \ALT_INV_Selector23~6_combout\,
	dataf => \ALT_INV_Equal3~11_combout\,
	combout => \Equal3~7_combout\);

-- Location: FF_X80_Y3_N13
\R.statusReg[0]_OTERM11_OTERM377_NEW_REG594\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Equal3~7_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.statusReg[0]_OTERM11_OTERM377_OTERM595\);

-- Location: FF_X80_Y6_N7
\R.statusReg[0]_OTERM11_OTERM377_NEW_REG592\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \vAluRes~52_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.statusReg[0]_OTERM11_OTERM377_OTERM593\);

-- Location: FF_X80_Y4_N26
\R.aluRes[24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Selector8~4_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(24));

-- Location: MLABCELL_X82_Y6_N6
\ShiftLeft0~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~29_combout\ = ( \R.aluData2\(2) & ( \ShiftLeft0~13_OTERM285\ & ( (!\R.aluData2\(3) & ((\ShiftLeft0~20_OTERM291\))) # (\R.aluData2\(3) & (\ShiftLeft0~8_OTERM207\)) ) ) ) # ( !\R.aluData2\(2) & ( \ShiftLeft0~13_OTERM285\ & ( (\R.aluData2\(3)) # 
-- (\ShiftLeft0~28_OTERM295\) ) ) ) # ( \R.aluData2\(2) & ( !\ShiftLeft0~13_OTERM285\ & ( (!\R.aluData2\(3) & ((\ShiftLeft0~20_OTERM291\))) # (\R.aluData2\(3) & (\ShiftLeft0~8_OTERM207\)) ) ) ) # ( !\R.aluData2\(2) & ( !\ShiftLeft0~13_OTERM285\ & ( 
-- (\ShiftLeft0~28_OTERM295\ & !\R.aluData2\(3)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100010001000100000000111100111101110111011101110000001111001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~28_OTERM295\,
	datab => \ALT_INV_R.aluData2\(3),
	datac => \ALT_INV_ShiftLeft0~8_OTERM207\,
	datad => \ALT_INV_ShiftLeft0~20_OTERM291\,
	datae => \ALT_INV_R.aluData2\(2),
	dataf => \ALT_INV_ShiftLeft0~13_OTERM285\,
	combout => \ShiftLeft0~29_combout\);

-- Location: LABCELL_X74_Y5_N6
\ShiftRight1~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~25_combout\ = ( \NxR.aluData2[0]~16_combout\ & ( \Mux236~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((\Mux235~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux233~0_combout\)) ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( 
-- \Mux236~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\) # (\Mux234~0_combout\) ) ) ) # ( \NxR.aluData2[0]~16_combout\ & ( !\Mux236~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((\Mux235~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & 
-- (\Mux233~0_combout\)) ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( !\Mux236~0_combout\ & ( (\Mux234~0_combout\ & \NxR.aluData2[1]~17_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000001011111010111110011111100110000010111110101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux233~0_combout\,
	datab => \ALT_INV_Mux234~0_combout\,
	datac => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datad => \ALT_INV_Mux235~0_combout\,
	datae => \ALT_INV_NxR.aluData2[0]~16_combout\,
	dataf => \ALT_INV_Mux236~0_combout\,
	combout => \ShiftRight1~25_combout\);

-- Location: FF_X74_Y5_N7
\ShiftRight1~25_NEW_REG276\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~25_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~25_OTERM277\);

-- Location: MLABCELL_X82_Y6_N24
\ShiftRight0~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight0~3_combout\ = ( \R.aluData2\(3) & ( \ShiftRight0~2_OTERM25\ & ( (\ShiftRight1~27_OTERM19\) # (\R.aluData2\(2)) ) ) ) # ( !\R.aluData2\(3) & ( \ShiftRight0~2_OTERM25\ & ( (!\R.aluData2\(2) & ((\ShiftRight1~25_OTERM277\))) # (\R.aluData2\(2) & 
-- (\ShiftRight1~26_OTERM37\)) ) ) ) # ( \R.aluData2\(3) & ( !\ShiftRight0~2_OTERM25\ & ( (!\R.aluData2\(2) & \ShiftRight1~27_OTERM19\) ) ) ) # ( !\R.aluData2\(3) & ( !\ShiftRight0~2_OTERM25\ & ( (!\R.aluData2\(2) & ((\ShiftRight1~25_OTERM277\))) # 
-- (\R.aluData2\(2) & (\ShiftRight1~26_OTERM37\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010110101111001000100010001000000101101011110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(2),
	datab => \ALT_INV_ShiftRight1~27_OTERM19\,
	datac => \ALT_INV_ShiftRight1~26_OTERM37\,
	datad => \ALT_INV_ShiftRight1~25_OTERM277\,
	datae => \ALT_INV_R.aluData2\(3),
	dataf => \ALT_INV_ShiftRight0~2_OTERM25\,
	combout => \ShiftRight0~3_combout\);

-- Location: MLABCELL_X82_Y6_N0
\Selector14~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector14~0_combout\ = ( \ShiftRight1~29_combout\ & ( \ShiftRight0~3_combout\ & ( (!\R.aluOp.ALUOpSRL~q\ & (!\R.aluOp.ALUOpSRA~q\ & ((!\R.aluOp.ALUOpSLL~q\) # (!\ShiftLeft0~29_combout\)))) ) ) ) # ( !\ShiftRight1~29_combout\ & ( \ShiftRight0~3_combout\ 
-- & ( (!\R.aluOp.ALUOpSRL~q\ & ((!\R.aluOp.ALUOpSLL~q\) # (!\ShiftLeft0~29_combout\))) ) ) ) # ( \ShiftRight1~29_combout\ & ( !\ShiftRight0~3_combout\ & ( (!\R.aluOp.ALUOpSRA~q\ & ((!\R.aluOp.ALUOpSLL~q\) # (!\ShiftLeft0~29_combout\))) ) ) ) # ( 
-- !\ShiftRight1~29_combout\ & ( !\ShiftRight0~3_combout\ & ( (!\R.aluOp.ALUOpSLL~q\) # (!\ShiftLeft0~29_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111110000110011001100000010101010101000001000100010000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpSRL~q\,
	datab => \ALT_INV_R.aluOp.ALUOpSRA~q\,
	datac => \ALT_INV_R.aluOp.ALUOpSLL~q\,
	datad => \ALT_INV_ShiftLeft0~29_combout\,
	datae => \ALT_INV_ShiftRight1~29_combout\,
	dataf => \ALT_INV_ShiftRight0~3_combout\,
	combout => \Selector14~0_combout\);

-- Location: LABCELL_X79_Y3_N6
\Selector14~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector14~5_combout\ = ( \Selector14~3_combout\ & ( (!\R.aluData2\(4) & !\Selector14~0_combout\) ) ) # ( !\Selector14~3_combout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111111111111111111111110000000000001111000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluData2\(4),
	datad => \ALT_INV_Selector14~0_combout\,
	dataf => \ALT_INV_Selector14~3_combout\,
	combout => \Selector14~5_combout\);

-- Location: FF_X79_Y3_N7
\R.aluRes[18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector14~5_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(18));

-- Location: FF_X80_Y4_N29
\R.aluRes[23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Selector9~5_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(23));

-- Location: LABCELL_X80_Y4_N51
\Selector14~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector14~4_combout\ = (!\Selector14~0_combout\ & !\R.aluData2\(4))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010000010100000101000001010000010100000101000001010000010100000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector14~0_combout\,
	datac => \ALT_INV_R.aluData2\(4),
	combout => \Selector14~4_combout\);

-- Location: LABCELL_X80_Y4_N45
\Equal3~12_RESYN1054\ : cyclonev_lcell_comb
-- Equation(s):
-- \Equal3~12_RESYN1054_BDD1055\ = ( \Selector14~4_combout\ & ( (!\R.aluRes\(24) & (!\R.aluCalc~q\ & (!\R.aluRes\(18) & !\R.aluRes\(23)))) ) ) # ( !\Selector14~4_combout\ & ( ((!\R.aluRes\(24) & (!\R.aluRes\(18) & !\R.aluRes\(23)))) # (\R.aluCalc~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1011001100110011101100110011001110000000000000001000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluRes\(24),
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_R.aluRes\(18),
	datad => \ALT_INV_R.aluRes\(23),
	dataf => \ALT_INV_Selector14~4_combout\,
	combout => \Equal3~12_RESYN1054_BDD1055\);

-- Location: LABCELL_X80_Y8_N6
\Equal3~12\ : cyclonev_lcell_comb
-- Equation(s):
-- \Equal3~12_combout\ = ( !\vAluRes~3_combout\ & ( !\vAluRes~5_combout\ & ( (!\vAluRes~10_combout\ & (!\vAluRes~4_combout\ & (\Equal3~12_RESYN1054_BDD1055\ & !\vAluRes~6_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000100000000000000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluRes~10_combout\,
	datab => \ALT_INV_vAluRes~4_combout\,
	datac => \ALT_INV_Equal3~12_RESYN1054_BDD1055\,
	datad => \ALT_INV_vAluRes~6_combout\,
	datae => \ALT_INV_vAluRes~3_combout\,
	dataf => \ALT_INV_vAluRes~5_combout\,
	combout => \Equal3~12_combout\);

-- Location: FF_X80_Y8_N7
\R.statusReg[0]_OTERM11_OTERM377_NEW_REG596\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Equal3~12_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.statusReg[0]_OTERM11_OTERM377_OTERM597\);

-- Location: LABCELL_X85_Y6_N12
\Equal3~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Equal3~13_combout\ = ( !\R.statusReg[0]_OTERM11_OTERM377_OTERM593\ & ( \R.statusReg[0]_OTERM11_OTERM377_OTERM597\ & ( \R.statusReg[0]_OTERM11_OTERM377_OTERM595\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000001111000011110000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.statusReg[0]_OTERM11_OTERM377_OTERM595\,
	datae => \ALT_INV_R.statusReg[0]_OTERM11_OTERM377_OTERM593\,
	dataf => \ALT_INV_R.statusReg[0]_OTERM11_OTERM377_OTERM597\,
	combout => \Equal3~13_combout\);

-- Location: MLABCELL_X84_Y4_N0
\Equal3~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Equal3~9_combout\ = ( \R.statusReg[0]_OTERM11_OTERM367\ & ( \Equal3~13_combout\ & ( (\R.statusReg[0]_OTERM11_OTERM375\ & (!\R.statusReg[0]_OTERM11_OTERM371\ & (\R.statusReg[0]_OTERM11_OTERM369\ & !\R.statusReg[0]_OTERM11_OTERM373\))) ) ) ) # ( 
-- !\R.statusReg[0]_OTERM11_OTERM367\ & ( \Equal3~13_combout\ & ( \R.statusReg[0]_OTERM11_OTERM375\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000001010101010101010000010000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.statusReg[0]_OTERM11_OTERM375\,
	datab => \ALT_INV_R.statusReg[0]_OTERM11_OTERM371\,
	datac => \ALT_INV_R.statusReg[0]_OTERM11_OTERM369\,
	datad => \ALT_INV_R.statusReg[0]_OTERM11_OTERM373\,
	datae => \ALT_INV_R.statusReg[0]_OTERM11_OTERM367\,
	dataf => \ALT_INV_Equal3~13_combout\,
	combout => \Equal3~9_combout\);

-- Location: FF_X77_Y3_N23
\R.aluRes[30]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector2~3_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes[30]~DUPLICATE_q\);

-- Location: LABCELL_X77_Y3_N48
\vAluRes~40\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~40_combout\ = ( !\R.aluCalc~q\ & ( (((\R.aluRes[30]~DUPLICATE_q\))) ) ) # ( \R.aluCalc~q\ & ( ((!\R.aluOp.ALUOpSub~q\ & (\R.aluOp.ALUOpAdd~q\ & (\Add1~121_sumout\))) # (\R.aluOp.ALUOpSub~q\ & (((\R.aluOp.ALUOpAdd~q\ & \Add1~121_sumout\)) # 
-- (\Add2~121_sumout\)))) # (\Selector2~2_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100001111010101010101111100001111000011110111011101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector2~2_combout\,
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_Add1~121_sumout\,
	datae => \ALT_INV_R.aluCalc~q\,
	dataf => \ALT_INV_Add2~121_sumout\,
	datag => \ALT_INV_R.aluRes[30]~DUPLICATE_q\,
	combout => \vAluRes~40_combout\);

-- Location: FF_X77_Y3_N49
\R.statusReg[0]_NEW_REG0\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \vAluRes~40_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.statusReg[0]_OTERM1\);

-- Location: LABCELL_X79_Y5_N27
\Add2~117\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~117_sumout\ = SUM(( !\R.aluData1\(29) $ (\R.aluData2\(29)) ) + ( \Add2~115\ ) + ( \Add2~114\ ))
-- \Add2~118\ = CARRY(( !\R.aluData1\(29) $ (\R.aluData2\(29)) ) + ( \Add2~115\ ) + ( \Add2~114\ ))
-- \Add2~119\ = SHARE((\R.aluData1\(29) & !\R.aluData2\(29)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010101010000000000000000000000001010101001010101",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData1\(29),
	datad => \ALT_INV_R.aluData2\(29),
	cin => \Add2~114\,
	sharein => \Add2~115\,
	sumout => \Add2~117_sumout\,
	cout => \Add2~118\,
	shareout => \Add2~119\);

-- Location: MLABCELL_X82_Y4_N54
\vAluRes~44\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~44_combout\ = ( !\R.aluCalc~q\ & ( (((\R.aluRes\(29)))) ) ) # ( \R.aluCalc~q\ & ( ((!\Add1~117_sumout\ & (\R.aluOp.ALUOpSub~q\ & ((\Add2~117_sumout\)))) # (\Add1~117_sumout\ & (((\R.aluOp.ALUOpSub~q\ & \Add2~117_sumout\)) # 
-- (\R.aluOp.ALUOpAdd~q\)))) # (\Selector3~2_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100001111000001011111111100001111000011110011011111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add1~117_sumout\,
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_Selector3~2_combout\,
	datae => \ALT_INV_R.aluCalc~q\,
	dataf => \ALT_INV_Add2~117_sumout\,
	datag => \ALT_INV_R.aluRes\(29),
	combout => \vAluRes~44_combout\);

-- Location: FF_X82_Y4_N56
\R.statusReg[0]_NEW_REG2\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \vAluRes~44_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.statusReg[0]_OTERM3\);

-- Location: LABCELL_X79_Y4_N48
\Equal3~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \Equal3~8_combout\ = ( !\R.statusReg[0]_OTERM1\ & ( !\R.statusReg[0]_OTERM3\ & ( (\Equal3~6_combout\ & (!\R.statusReg[0]_OTERM5\ & (\Equal3~2_combout\ & \Equal3~9_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000100000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Equal3~6_combout\,
	datab => \ALT_INV_R.statusReg[0]_OTERM5\,
	datac => \ALT_INV_Equal3~2_combout\,
	datad => \ALT_INV_Equal3~9_combout\,
	datae => \ALT_INV_R.statusReg[0]_OTERM1\,
	dataf => \ALT_INV_R.statusReg[0]_OTERM3\,
	combout => \Equal3~8_combout\);

-- Location: LABCELL_X79_Y4_N30
\vAluRes~36\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~36_combout\ = ( !\R.aluCalc~q\ & ( (((\R.aluRes\(31)))) ) ) # ( \R.aluCalc~q\ & ( ((!\R.aluOp.ALUOpSub~q\ & (((\R.aluOp.ALUOpAdd~q\ & \Add1~125_sumout\)))) # (\R.aluOp.ALUOpSub~q\ & (((\R.aluOp.ALUOpAdd~q\ & \Add1~125_sumout\)) # 
-- (\Add2~125_sumout\)))) # (\Selector1~2_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100001111000100011111111100001111000011110001111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datab => \ALT_INV_Add2~125_sumout\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_Selector1~2_combout\,
	datae => \ALT_INV_R.aluCalc~q\,
	dataf => \ALT_INV_Add1~125_sumout\,
	datag => \ALT_INV_R.aluRes\(31),
	combout => \vAluRes~36_combout\);

-- Location: FF_X79_Y4_N32
\R.statusReg[1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \vAluRes~36_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.statusReg\(1));

-- Location: LABCELL_X81_Y7_N42
\ShiftLeft0~57\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~57_combout\ = ( \R.aluData2\(1) & ( \R.aluData1\(29) & ( (\R.aluData1\(30)) # (\R.aluData2\(0)) ) ) ) # ( !\R.aluData2\(1) & ( \R.aluData1\(29) & ( (\R.aluData1\(31) & \R.aluData2\(0)) ) ) ) # ( \R.aluData2\(1) & ( !\R.aluData1\(29) & ( 
-- (!\R.aluData2\(0) & \R.aluData1\(30)) ) ) ) # ( !\R.aluData2\(1) & ( !\R.aluData1\(29) & ( (\R.aluData1\(31) & \R.aluData2\(0)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100010001000011000000110000010001000100010011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData1\(31),
	datab => \ALT_INV_R.aluData2\(0),
	datac => \ALT_INV_R.aluData1\(30),
	datae => \ALT_INV_R.aluData2\(1),
	dataf => \ALT_INV_R.aluData1\(29),
	combout => \ShiftLeft0~57_combout\);

-- Location: LABCELL_X81_Y8_N0
\ShiftLeft0~58\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~58_combout\ = ( \ShiftLeft0~49_OTERM761\ & ( \ShiftLeft0~57_combout\ & ( (!\R.aluData2\(3)) # ((!\R.aluData2\(2) & ((\ShiftLeft0~40_OTERM755\))) # (\R.aluData2\(2) & (\ShiftLeft0~32_OTERM297\))) ) ) ) # ( !\ShiftLeft0~49_OTERM761\ & ( 
-- \ShiftLeft0~57_combout\ & ( (!\R.aluData2\(2) & (((!\R.aluData2\(3)) # (\ShiftLeft0~40_OTERM755\)))) # (\R.aluData2\(2) & (\ShiftLeft0~32_OTERM297\ & (\R.aluData2\(3)))) ) ) ) # ( \ShiftLeft0~49_OTERM761\ & ( !\ShiftLeft0~57_combout\ & ( (!\R.aluData2\(2) 
-- & (((\R.aluData2\(3) & \ShiftLeft0~40_OTERM755\)))) # (\R.aluData2\(2) & (((!\R.aluData2\(3))) # (\ShiftLeft0~32_OTERM297\))) ) ) ) # ( !\ShiftLeft0~49_OTERM761\ & ( !\ShiftLeft0~57_combout\ & ( (\R.aluData2\(3) & ((!\R.aluData2\(2) & 
-- ((\ShiftLeft0~40_OTERM755\))) # (\R.aluData2\(2) & (\ShiftLeft0~32_OTERM297\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000100001011010100010101101110100001101010111111000111111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(2),
	datab => \ALT_INV_ShiftLeft0~32_OTERM297\,
	datac => \ALT_INV_R.aluData2\(3),
	datad => \ALT_INV_ShiftLeft0~40_OTERM755\,
	datae => \ALT_INV_ShiftLeft0~49_OTERM761\,
	dataf => \ALT_INV_ShiftLeft0~57_combout\,
	combout => \ShiftLeft0~58_combout\);

-- Location: LABCELL_X81_Y8_N6
\Selector0~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector0~0_combout\ = ( \ShiftLeft0~58_combout\ & ( \R.aluData1\(31) & ( ((\R.aluOp.ALUOpSLL~q\ & ((!\R.aluData2\(4)) # (\ShiftLeft0~25_combout\)))) # (\R.aluOp.ALUOpSRA~q\) ) ) ) # ( !\ShiftLeft0~58_combout\ & ( \R.aluData1\(31) & ( ((\R.aluData2\(4) & 
-- (\ShiftLeft0~25_combout\ & \R.aluOp.ALUOpSLL~q\))) # (\R.aluOp.ALUOpSRA~q\) ) ) ) # ( \ShiftLeft0~58_combout\ & ( !\R.aluData1\(31) & ( (\R.aluOp.ALUOpSLL~q\ & ((!\R.aluData2\(4)) # (\ShiftLeft0~25_combout\))) ) ) ) # ( !\ShiftLeft0~58_combout\ & ( 
-- !\R.aluData1\(31) & ( (\R.aluData2\(4) & (\ShiftLeft0~25_combout\ & \R.aluOp.ALUOpSLL~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000101000000001010111100110011001101110011001110111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(4),
	datab => \ALT_INV_R.aluOp.ALUOpSRA~q\,
	datac => \ALT_INV_ShiftLeft0~25_combout\,
	datad => \ALT_INV_R.aluOp.ALUOpSLL~q\,
	datae => \ALT_INV_ShiftLeft0~58_combout\,
	dataf => \ALT_INV_R.aluData1\(31),
	combout => \Selector0~0_combout\);

-- Location: MLABCELL_X78_Y5_N36
\Add1~129\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~129_sumout\ = SUM(( GND ) + ( GND ) + ( \Add1~126\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	cin => \Add1~126\,
	sumout => \Add1~129_sumout\);

-- Location: LABCELL_X79_Y5_N30
\Add2~121\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~121_sumout\ = SUM(( !\R.aluData1\(30) $ (\R.aluData2\(30)) ) + ( \Add2~119\ ) + ( \Add2~118\ ))
-- \Add2~122\ = CARRY(( !\R.aluData1\(30) $ (\R.aluData2\(30)) ) + ( \Add2~119\ ) + ( \Add2~118\ ))
-- \Add2~123\ = SHARE((\R.aluData1\(30) & !\R.aluData2\(30)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000001100110000000000000000000000001100110000110011",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluData1\(30),
	datad => \ALT_INV_R.aluData2\(30),
	cin => \Add2~118\,
	sharein => \Add2~119\,
	sumout => \Add2~121_sumout\,
	cout => \Add2~122\,
	shareout => \Add2~123\);

-- Location: LABCELL_X79_Y5_N33
\Add2~125\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~125_sumout\ = SUM(( !\R.aluData2\(31) $ (\R.aluData1\(31)) ) + ( \Add2~123\ ) + ( \Add2~122\ ))
-- \Add2~126\ = CARRY(( !\R.aluData2\(31) $ (\R.aluData1\(31)) ) + ( \Add2~123\ ) + ( \Add2~122\ ))
-- \Add2~127\ = SHARE((!\R.aluData2\(31) & \R.aluData1\(31)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000001111000000000000000000001111000000001111",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluData2\(31),
	datad => \ALT_INV_R.aluData1\(31),
	cin => \Add2~122\,
	sharein => \Add2~123\,
	sumout => \Add2~125_sumout\,
	cout => \Add2~126\,
	shareout => \Add2~127\);

-- Location: LABCELL_X79_Y5_N36
\Add2~129\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add2~129_sumout\ = SUM(( VCC ) + ( \Add2~127\ ) + ( \Add2~126\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000001111111111111111",
	shared_arith => "on")
-- pragma translate_on
PORT MAP (
	cin => \Add2~126\,
	sharein => \Add2~127\,
	sumout => \Add2~129_sumout\);

-- Location: LABCELL_X79_Y4_N54
\Selector0~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector0~1_combout\ = ( \Add1~129_sumout\ & ( \Add2~129_sumout\ & ( ((\Selector0~0_combout\) # (\R.aluOp.ALUOpSub~q\)) # (\R.aluOp.ALUOpAdd~q\) ) ) ) # ( !\Add1~129_sumout\ & ( \Add2~129_sumout\ & ( (\Selector0~0_combout\) # (\R.aluOp.ALUOpSub~q\) ) ) ) 
-- # ( \Add1~129_sumout\ & ( !\Add2~129_sumout\ & ( (\Selector0~0_combout\) # (\R.aluOp.ALUOpAdd~q\) ) ) ) # ( !\Add1~129_sumout\ & ( !\Add2~129_sumout\ & ( \Selector0~0_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111010101011111111100001111111111110101111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datac => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datad => \ALT_INV_Selector0~0_combout\,
	datae => \ALT_INV_Add1~129_sumout\,
	dataf => \ALT_INV_Add2~129_sumout\,
	combout => \Selector0~1_combout\);

-- Location: FF_X79_Y4_N56
\R.statusReg[2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector0~1_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.statusReg\(2));

-- Location: LABCELL_X79_Y4_N24
\Mux58~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux58~0_combout\ = ( \R.statusReg\(2) & ( \R.curInst\(13) & ( (\R.curInst\(14) & !\R.curInst\(12)) ) ) ) # ( !\R.statusReg\(2) & ( \R.curInst\(13) & ( (\R.curInst\(14) & \R.curInst\(12)) ) ) ) # ( \R.statusReg\(2) & ( !\R.curInst\(13) & ( 
-- !\R.curInst\(12) $ (((!\R.curInst\(14) & (!\Equal3~8_combout\)) # (\R.curInst\(14) & ((!\R.statusReg\(1)))))) ) ) ) # ( !\R.statusReg\(2) & ( !\R.curInst\(13) & ( !\R.curInst\(12) $ (((!\R.curInst\(14) & (!\Equal3~8_combout\)) # (\R.curInst\(14) & 
-- ((!\R.statusReg\(1)))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100101101111000010010110111100000000011000000110011000000110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Equal3~8_combout\,
	datab => \ALT_INV_R.curInst\(14),
	datac => \ALT_INV_R.curInst\(12),
	datad => \ALT_INV_R.statusReg\(1),
	datae => \ALT_INV_R.statusReg\(2),
	dataf => \ALT_INV_R.curInst\(13),
	combout => \Mux58~0_combout\);

-- Location: LABCELL_X79_Y4_N36
\NxR~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR~8_combout\ = ( \Mux58~0_combout\ & ( (!\R.ctrlState.ReadReg~q\ & (\R.ctrlState.CheckJump~q\)) # (\R.ctrlState.ReadReg~q\ & (((\Equal4~0_combout\ & \Equal4~1_combout\)))) ) ) # ( !\Mux58~0_combout\ & ( (\R.ctrlState.ReadReg~q\ & (\Equal4~0_combout\ & 
-- \Equal4~1_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000101000000000000010100100010001001110010001000100111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.ctrlState.ReadReg~q\,
	datab => \ALT_INV_R.ctrlState.CheckJump~q\,
	datac => \ALT_INV_Equal4~0_combout\,
	datad => \ALT_INV_Equal4~1_combout\,
	dataf => \ALT_INV_Mux58~0_combout\,
	combout => \NxR~8_combout\);

-- Location: FF_X79_Y4_N38
\R.jumpToAdr\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR~8_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sclr => \R.ctrlState.Fetch~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.jumpToAdr~q\);

-- Location: FF_X82_Y7_N8
\R.regWriteData[5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \R.regWriteData[5]~feeder_combout\,
	asdata => \Comb:vRegWriteData[5]~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(5));

-- Location: FF_X60_Y7_N20
\RegFile[29][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(5),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][5]~q\);

-- Location: LABCELL_X62_Y7_N42
\Mux85~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux85~22_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & (\RegFile[24][5]~q\)) # (\R.curInst\(15) & ((\RegFile[25][5]~q\))))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & ((\RegFile[26][5]~q\))) # (\R.curInst\(15) & (\RegFile[27][5]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110000110011111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[27][5]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[26][5]~q\,
	datad => \ALT_INV_RegFile[25][5]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][5]~q\,
	combout => \Mux85~22_combout\);

-- Location: LABCELL_X62_Y7_N30
\Mux85~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux85~9_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux85~22_combout\)))) # (\R.curInst\(17) & ((!\Mux85~22_combout\ & ((\RegFile[28][5]~q\))) # (\Mux85~22_combout\ & (\RegFile[29][5]~q\))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) 
-- & (((\Mux85~22_combout\)))) # (\R.curInst\(17) & ((!\Mux85~22_combout\ & ((\RegFile[30][5]~q\))) # (\Mux85~22_combout\ & (\RegFile[31][5]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[29][5]~q\,
	datab => \ALT_INV_RegFile[31][5]~q\,
	datac => \ALT_INV_RegFile[30][5]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux85~22_combout\,
	datag => \ALT_INV_RegFile[28][5]~q\,
	combout => \Mux85~9_combout\);

-- Location: MLABCELL_X65_Y3_N36
\Mux85~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux85~14_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[8][5]~q\))) # (\R.curInst\(15) & (\RegFile[9][5]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[10][5]~q\))) # (\R.curInst\(15) & (\RegFile[11][5]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[11][5]~q\,
	datab => \ALT_INV_RegFile[9][5]~q\,
	datac => \ALT_INV_RegFile[10][5]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][5]~q\,
	combout => \Mux85~14_combout\);

-- Location: LABCELL_X66_Y7_N42
\Mux85~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux85~1_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux85~14_combout\)))) # (\R.curInst\(17) & ((!\Mux85~14_combout\ & ((\RegFile[12][5]~q\))) # (\Mux85~14_combout\ & (\RegFile[13][5]~q\))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) 
-- & (((\Mux85~14_combout\)))) # (\R.curInst\(17) & ((!\Mux85~14_combout\ & ((\RegFile[14][5]~q\))) # (\Mux85~14_combout\ & (\RegFile[15][5]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][5]~q\,
	datab => \ALT_INV_RegFile[13][5]~q\,
	datac => \ALT_INV_RegFile[14][5]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux85~14_combout\,
	datag => \ALT_INV_RegFile[12][5]~q\,
	combout => \Mux85~1_combout\);

-- Location: LABCELL_X62_Y7_N24
\Mux85~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux85~0_combout\ = ( \RegFile[4][5]~q\ & ( \R.curInst\(15) & ( (!\R.curInst\(16) & (\RegFile[5][5]~q\)) # (\R.curInst\(16) & ((\RegFile[7][5]~q\))) ) ) ) # ( !\RegFile[4][5]~q\ & ( \R.curInst\(15) & ( (!\R.curInst\(16) & (\RegFile[5][5]~q\)) # 
-- (\R.curInst\(16) & ((\RegFile[7][5]~q\))) ) ) ) # ( \RegFile[4][5]~q\ & ( !\R.curInst\(15) & ( (!\R.curInst\(16)) # (\RegFile[6][5]~q\) ) ) ) # ( !\RegFile[4][5]~q\ & ( !\R.curInst\(15) & ( (\RegFile[6][5]~q\ & \R.curInst\(16)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110011111111110011001101010101000011110101010100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[5][5]~q\,
	datab => \ALT_INV_RegFile[6][5]~q\,
	datac => \ALT_INV_RegFile[7][5]~q\,
	datad => \ALT_INV_R.curInst\(16),
	datae => \ALT_INV_RegFile[4][5]~q\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux85~0_combout\);

-- Location: LABCELL_X62_Y7_N12
\Mux85~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux85~26_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (\R.curInst\(15) & (\RegFile[1][5]~q\))) # (\R.curInst\(17) & ((((\Mux85~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & ((!\R.curInst\(15) & (\RegFile[2][5]~q\)) # 
-- (\R.curInst\(15) & (((\RegFile[3][5]~q\)))))) # (\R.curInst\(17) & ((((\Mux85~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010000000100000010000100110000110111001101110011101101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(15),
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[2][5]~q\,
	datad => \ALT_INV_RegFile[3][5]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux85~0_combout\,
	datag => \ALT_INV_RegFile[1][5]~q\,
	combout => \Mux85~26_combout\);

-- Location: FF_X60_Y7_N56
\RegFile[16][5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[16][5]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][5]~q\);

-- Location: LABCELL_X63_Y7_N30
\Mux85~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux85~18_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[16][5]~q\))) # (\R.curInst\(15) & (\RegFile[17][5]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[18][5]~q\))) # (\R.curInst\(15) & (\RegFile[19][5]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[17][5]~q\,
	datab => \ALT_INV_RegFile[19][5]~q\,
	datac => \ALT_INV_RegFile[18][5]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][5]~q\,
	combout => \Mux85~18_combout\);

-- Location: LABCELL_X63_Y7_N27
\Mux85~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux85~5_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux85~18_combout\))))) # (\R.curInst\(17) & (((!\Mux85~18_combout\ & (\RegFile[20][5]~q\)) # (\Mux85~18_combout\ & ((\RegFile[21][5]~q\)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) 
-- & ((((\Mux85~18_combout\))))) # (\R.curInst\(17) & (((!\Mux85~18_combout\ & ((\RegFile[22][5]~q\))) # (\Mux85~18_combout\ & (\RegFile[23][5]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110101010111111111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[23][5]~q\,
	datac => \ALT_INV_RegFile[22][5]~q\,
	datad => \ALT_INV_RegFile[21][5]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux85~18_combout\,
	datag => \ALT_INV_RegFile[20][5]~q\,
	combout => \Mux85~5_combout\);

-- Location: LABCELL_X66_Y7_N54
\Mux85~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux85~13_combout\ = ( \Mux85~26_combout\ & ( \Mux85~5_combout\ & ( (!\R.curInst\(18)) # ((!\R.curInst\(19) & ((\Mux85~1_combout\))) # (\R.curInst\(19) & (\Mux85~9_combout\))) ) ) ) # ( !\Mux85~26_combout\ & ( \Mux85~5_combout\ & ( (!\R.curInst\(18) & 
-- (((\R.curInst\(19))))) # (\R.curInst\(18) & ((!\R.curInst\(19) & ((\Mux85~1_combout\))) # (\R.curInst\(19) & (\Mux85~9_combout\)))) ) ) ) # ( \Mux85~26_combout\ & ( !\Mux85~5_combout\ & ( (!\R.curInst\(18) & (((!\R.curInst\(19))))) # (\R.curInst\(18) & 
-- ((!\R.curInst\(19) & ((\Mux85~1_combout\))) # (\R.curInst\(19) & (\Mux85~9_combout\)))) ) ) ) # ( !\Mux85~26_combout\ & ( !\Mux85~5_combout\ & ( (\R.curInst\(18) & ((!\R.curInst\(19) & ((\Mux85~1_combout\))) # (\R.curInst\(19) & (\Mux85~9_combout\)))) ) ) 
-- )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000101010001101000011111000100001011010110111010101111111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(18),
	datab => \ALT_INV_Mux85~9_combout\,
	datac => \ALT_INV_R.curInst\(19),
	datad => \ALT_INV_Mux85~1_combout\,
	datae => \ALT_INV_Mux85~26_combout\,
	dataf => \ALT_INV_Mux85~5_combout\,
	combout => \Mux85~13_combout\);

-- Location: LABCELL_X73_Y7_N51
\Mux249~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux249~0_combout\ = ( !\vAluSrc1~1_combout\ & ( \Mux85~13_combout\ & ( (!\vAluSrc1~2_combout\) # (\R.curPC\(5)) ) ) ) # ( !\vAluSrc1~1_combout\ & ( !\Mux85~13_combout\ & ( (\R.curPC\(5) & \vAluSrc1~2_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000000000000011110011111100110000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.curPC\(5),
	datac => \ALT_INV_vAluSrc1~2_combout\,
	datae => \ALT_INV_vAluSrc1~1_combout\,
	dataf => \ALT_INV_Mux85~13_combout\,
	combout => \Mux249~0_combout\);

-- Location: LABCELL_X73_Y7_N42
\ShiftLeft0~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~8_combout\ = ( \NxR.aluData2[0]~16_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( \Mux251~0_combout\ ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( \Mux250~0_combout\ ) ) ) # ( \NxR.aluData2[0]~16_combout\ & ( 
-- !\NxR.aluData2[1]~17_combout\ & ( \Mux249~0_combout\ ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( !\NxR.aluData2[1]~17_combout\ & ( \Mux248~0_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101000000001111111100110011001100110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux248~0_combout\,
	datab => \ALT_INV_Mux250~0_combout\,
	datac => \ALT_INV_Mux251~0_combout\,
	datad => \ALT_INV_Mux249~0_combout\,
	datae => \ALT_INV_NxR.aluData2[0]~16_combout\,
	dataf => \ALT_INV_NxR.aluData2[1]~17_combout\,
	combout => \ShiftLeft0~8_combout\);

-- Location: FF_X73_Y7_N43
\ShiftLeft0~8_NEW_REG206\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~8_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~8_OTERM207\);

-- Location: MLABCELL_X82_Y6_N15
\Selector26~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector26~1_combout\ = ( \ShiftLeft0~8_OTERM207\ & ( (!\R.aluData2\(3) & (\Selector27~0_OTERM385\ & ((!\R.aluData2\(2)) # (\ShiftLeft0~2_OTERM221\)))) ) ) # ( !\ShiftLeft0~8_OTERM207\ & ( (\R.aluData2\(2) & (!\R.aluData2\(3) & (\ShiftLeft0~2_OTERM221\ & 
-- \Selector27~0_OTERM385\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000100000000000000010000000000100011000000000010001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(2),
	datab => \ALT_INV_R.aluData2\(3),
	datac => \ALT_INV_ShiftLeft0~2_OTERM221\,
	datad => \ALT_INV_Selector27~0_OTERM385\,
	dataf => \ALT_INV_ShiftLeft0~8_OTERM207\,
	combout => \Selector26~1_combout\);

-- Location: MLABCELL_X82_Y6_N12
\ShiftRight0~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight0~9_combout\ = ( \ShiftRight1~27_OTERM19\ & ( (!\R.aluData2\(2) & ((!\R.aluData2\(3) & (\ShiftRight1~26_OTERM37\)) # (\R.aluData2\(3) & ((\ShiftRight0~2_OTERM25\))))) # (\R.aluData2\(2) & (!\R.aluData2\(3))) ) ) # ( !\ShiftRight1~27_OTERM19\ & 
-- ( (!\R.aluData2\(2) & ((!\R.aluData2\(3) & (\ShiftRight1~26_OTERM37\)) # (\R.aluData2\(3) & ((\ShiftRight0~2_OTERM25\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000100000101010000010000010101001001100011011100100110001101110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(2),
	datab => \ALT_INV_R.aluData2\(3),
	datac => \ALT_INV_ShiftRight1~26_OTERM37\,
	datad => \ALT_INV_ShiftRight0~2_OTERM25\,
	dataf => \ALT_INV_ShiftRight1~27_OTERM19\,
	combout => \ShiftRight0~9_combout\);

-- Location: LABCELL_X74_Y6_N48
\ShiftRight1~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~22_combout\ = ( \Mux243~0_combout\ & ( \Mux244~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\) # ((!\NxR.aluData2[0]~16_combout\ & ((\Mux242~0_combout\))) # (\NxR.aluData2[0]~16_combout\ & (\Mux241~0_combout\))) ) ) ) # ( !\Mux243~0_combout\ & 
-- ( \Mux244~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((!\NxR.aluData2[0]~16_combout\)))) # (\NxR.aluData2[1]~17_combout\ & ((!\NxR.aluData2[0]~16_combout\ & ((\Mux242~0_combout\))) # (\NxR.aluData2[0]~16_combout\ & (\Mux241~0_combout\)))) ) ) ) # ( 
-- \Mux243~0_combout\ & ( !\Mux244~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((\NxR.aluData2[0]~16_combout\)))) # (\NxR.aluData2[1]~17_combout\ & ((!\NxR.aluData2[0]~16_combout\ & ((\Mux242~0_combout\))) # (\NxR.aluData2[0]~16_combout\ & 
-- (\Mux241~0_combout\)))) ) ) ) # ( !\Mux243~0_combout\ & ( !\Mux244~0_combout\ & ( (\NxR.aluData2[1]~17_combout\ & ((!\NxR.aluData2[0]~16_combout\ & ((\Mux242~0_combout\))) # (\NxR.aluData2[0]~16_combout\ & (\Mux241~0_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100010001000001011011101110101111000100011010111110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datab => \ALT_INV_Mux241~0_combout\,
	datac => \ALT_INV_Mux242~0_combout\,
	datad => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datae => \ALT_INV_Mux243~0_combout\,
	dataf => \ALT_INV_Mux244~0_combout\,
	combout => \ShiftRight1~22_combout\);

-- Location: FF_X74_Y6_N49
\ShiftRight1~22_NEW_REG272\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~22_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~22_OTERM273\);

-- Location: LABCELL_X73_Y6_N51
\ShiftRight1~23\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~23_combout\ = ( \Mux238~0_combout\ & ( \NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((\Mux239~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux237~0_combout\)) ) ) ) # ( !\Mux238~0_combout\ & ( 
-- \NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((\Mux239~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux237~0_combout\)) ) ) ) # ( \Mux238~0_combout\ & ( !\NxR.aluData2[0]~16_combout\ & ( (\NxR.aluData2[1]~17_combout\) # 
-- (\Mux240~0_combout\) ) ) ) # ( !\Mux238~0_combout\ & ( !\NxR.aluData2[0]~16_combout\ & ( (\Mux240~0_combout\ & !\NxR.aluData2[1]~17_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100000000001100111111111100001111010101010000111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux237~0_combout\,
	datab => \ALT_INV_Mux240~0_combout\,
	datac => \ALT_INV_Mux239~0_combout\,
	datad => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datae => \ALT_INV_Mux238~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[0]~16_combout\,
	combout => \ShiftRight1~23_combout\);

-- Location: FF_X73_Y6_N53
\ShiftRight1~23_NEW_REG274\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~23_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~23_OTERM275\);

-- Location: LABCELL_X75_Y7_N36
\ShiftRight1~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~21_combout\ = ( \Mux245~0_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( (\NxR.aluData2[0]~16_combout\) # (\Mux246~0_combout\) ) ) ) # ( !\Mux245~0_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( (\Mux246~0_combout\ & 
-- !\NxR.aluData2[0]~16_combout\) ) ) ) # ( \Mux245~0_combout\ & ( !\NxR.aluData2[1]~17_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (\Mux248~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & ((\Mux247~0_combout\))) ) ) ) # ( !\Mux245~0_combout\ & ( 
-- !\NxR.aluData2[1]~17_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (\Mux248~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & ((\Mux247~0_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010100110011010101010011001100001111000000000000111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux248~0_combout\,
	datab => \ALT_INV_Mux247~0_combout\,
	datac => \ALT_INV_Mux246~0_combout\,
	datad => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datae => \ALT_INV_Mux245~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[1]~17_combout\,
	combout => \ShiftRight1~21_combout\);

-- Location: FF_X75_Y7_N37
\ShiftRight1~21_NEW_REG270\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~21_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~21_OTERM271\);

-- Location: MLABCELL_X84_Y6_N36
\ShiftRight1~44\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~44_combout\ = ( \ShiftRight1~25_OTERM277\ & ( \ShiftRight1~21_OTERM271\ & ( (!\R.aluData2\(3) & (((!\R.aluData2\(2))) # (\ShiftRight1~22_OTERM273\))) # (\R.aluData2\(3) & (((\R.aluData2\(2)) # (\ShiftRight1~23_OTERM275\)))) ) ) ) # ( 
-- !\ShiftRight1~25_OTERM277\ & ( \ShiftRight1~21_OTERM271\ & ( (!\R.aluData2\(3) & (((!\R.aluData2\(2))) # (\ShiftRight1~22_OTERM273\))) # (\R.aluData2\(3) & (((\ShiftRight1~23_OTERM275\ & !\R.aluData2\(2))))) ) ) ) # ( \ShiftRight1~25_OTERM277\ & ( 
-- !\ShiftRight1~21_OTERM271\ & ( (!\R.aluData2\(3) & (\ShiftRight1~22_OTERM273\ & ((\R.aluData2\(2))))) # (\R.aluData2\(3) & (((\R.aluData2\(2)) # (\ShiftRight1~23_OTERM275\)))) ) ) ) # ( !\ShiftRight1~25_OTERM277\ & ( !\ShiftRight1~21_OTERM271\ & ( 
-- (!\R.aluData2\(3) & (\ShiftRight1~22_OTERM273\ & ((\R.aluData2\(2))))) # (\R.aluData2\(3) & (((\ShiftRight1~23_OTERM275\ & !\R.aluData2\(2))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100100010000001010111011110101111001000101010111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(3),
	datab => \ALT_INV_ShiftRight1~22_OTERM273\,
	datac => \ALT_INV_ShiftRight1~23_OTERM275\,
	datad => \ALT_INV_R.aluData2\(2),
	datae => \ALT_INV_ShiftRight1~25_OTERM277\,
	dataf => \ALT_INV_ShiftRight1~21_OTERM271\,
	combout => \ShiftRight1~44_combout\);

-- Location: MLABCELL_X82_Y6_N54
\Selector26~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector26~3_combout\ = ( !\Selector31~5_OTERM599\ & ( \ShiftRight1~44_combout\ & ( (!\Selector26~2_OTERM415\ & (!\Selector26~1_combout\ & ((!\Selector31~7_OTERM383\) # (!\ShiftRight0~9_combout\)))) ) ) ) # ( \Selector31~5_OTERM599\ & ( 
-- !\ShiftRight1~44_combout\ & ( (!\Selector26~2_OTERM415\ & (!\Selector26~1_combout\ & ((!\Selector31~7_OTERM383\) # (!\ShiftRight0~9_combout\)))) ) ) ) # ( !\Selector31~5_OTERM599\ & ( !\ShiftRight1~44_combout\ & ( (!\Selector26~2_OTERM415\ & 
-- (!\Selector26~1_combout\ & ((!\Selector31~7_OTERM383\) # (!\ShiftRight0~9_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000100010000000100010001000000010001000100000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector26~2_OTERM415\,
	datab => \ALT_INV_Selector26~1_combout\,
	datac => \ALT_INV_Selector31~7_OTERM383\,
	datad => \ALT_INV_ShiftRight0~9_combout\,
	datae => \ALT_INV_Selector31~5_OTERM599\,
	dataf => \ALT_INV_ShiftRight1~44_combout\,
	combout => \Selector26~3_combout\);

-- Location: MLABCELL_X78_Y6_N18
\Add1~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~25_sumout\ = SUM(( \Add2~25_OTERM723_OTERM833\ ) + ( \Add2~25_OTERM723_OTERM835\ ) + ( \Add1~22\ ))
-- \Add1~26\ = CARRY(( \Add2~25_OTERM723_OTERM833\ ) + ( \Add2~25_OTERM723_OTERM835\ ) + ( \Add1~22\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Add2~25_OTERM723_OTERM835\,
	datad => \ALT_INV_Add2~25_OTERM723_OTERM833\,
	cin => \Add1~22\,
	sumout => \Add1~25_sumout\,
	cout => \Add1~26\);

-- Location: LABCELL_X83_Y6_N6
\Selector26~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector26~0_combout\ = ( \Add1~25_sumout\ & ( ((\R.aluOp.ALUOpSub~q\ & \Add2~25_sumout\)) # (\R.aluOp.ALUOpAdd~q\) ) ) # ( !\Add1~25_sumout\ & ( (\R.aluOp.ALUOpSub~q\ & \Add2~25_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110011000000000011001100001111001111110000111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_Add2~25_sumout\,
	dataf => \ALT_INV_Add1~25_sumout\,
	combout => \Selector26~0_combout\);

-- Location: IOIBUF_X36_Y81_N35
\avm_d_readdata[30]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(30),
	o => \avm_d_readdata[30]~input_o\);

-- Location: LABCELL_X80_Y6_N21
\Comb:vRegWriteData[6]~0_RESYN1098\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[6]~0_RESYN1098_BDD1099\ = ( \ShiftRight1~43_combout\ & ( \R.aluRes\(6) & ( (!\R.memToReg~q\ & ((!\R.aluCalc~q\) # ((\Selector31~6_OTERM381\)))) # (\R.memToReg~q\ & (((\Mux222~0_combout\)))) ) ) ) # ( !\ShiftRight1~43_combout\ & ( 
-- \R.aluRes\(6) & ( (!\R.memToReg~q\ & (!\R.aluCalc~q\)) # (\R.memToReg~q\ & ((\Mux222~0_combout\))) ) ) ) # ( \ShiftRight1~43_combout\ & ( !\R.aluRes\(6) & ( (!\R.memToReg~q\ & (\R.aluCalc~q\ & ((\Selector31~6_OTERM381\)))) # (\R.memToReg~q\ & 
-- (((\Mux222~0_combout\)))) ) ) ) # ( !\ShiftRight1~43_combout\ & ( !\R.aluRes\(6) & ( (\Mux222~0_combout\ & \R.memToReg~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110011000001010011001110101010001100111010111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluCalc~q\,
	datab => \ALT_INV_Mux222~0_combout\,
	datac => \ALT_INV_Selector31~6_OTERM381\,
	datad => \ALT_INV_R.memToReg~q\,
	datae => \ALT_INV_ShiftRight1~43_combout\,
	dataf => \ALT_INV_R.aluRes\(6),
	combout => \Comb:vRegWriteData[6]~0_RESYN1098_BDD1099\);

-- Location: LABCELL_X83_Y6_N18
\Comb:vRegWriteData[6]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[6]~0_combout\ = ( \avm_d_readdata[30]~input_o\ & ( \Comb:vRegWriteData[6]~0_RESYN1098_BDD1099\ ) ) # ( !\avm_d_readdata[30]~input_o\ & ( \Comb:vRegWriteData[6]~0_RESYN1098_BDD1099\ & ( !\R.memToReg~q\ ) ) ) # ( 
-- \avm_d_readdata[30]~input_o\ & ( !\Comb:vRegWriteData[6]~0_RESYN1098_BDD1099\ & ( (!\R.memToReg~q\ & (\R.aluCalc~q\ & ((!\Selector26~3_combout\) # (\Selector26~0_combout\)))) ) ) ) # ( !\avm_d_readdata[30]~input_o\ & ( 
-- !\Comb:vRegWriteData[6]~0_RESYN1098_BDD1099\ & ( (!\R.memToReg~q\ & (\R.aluCalc~q\ & ((!\Selector26~3_combout\) # (\Selector26~0_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000100000001010000010000000101010101010101010101111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.memToReg~q\,
	datab => \ALT_INV_Selector26~3_combout\,
	datac => \ALT_INV_R.aluCalc~q\,
	datad => \ALT_INV_Selector26~0_combout\,
	datae => \ALT_INV_avm_d_readdata[30]~input_o\,
	dataf => \ALT_INV_Comb:vRegWriteData[6]~0_RESYN1098_BDD1099\,
	combout => \Comb:vRegWriteData[6]~0_combout\);

-- Location: FF_X83_Y6_N29
\R.regWriteData[6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \R.regWriteData[6]~feeder_combout\,
	asdata => \Comb:vRegWriteData[6]~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(6));

-- Location: FF_X65_Y8_N38
\RegFile[21][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(6),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][6]~q\);

-- Location: FF_X64_Y7_N32
\RegFile[23][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(6),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][6]~q\);

-- Location: FF_X64_Y4_N4
\RegFile[22][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(6),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][6]~q\);

-- Location: FF_X65_Y8_N20
\RegFile[17][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(6),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][6]~q\);

-- Location: LABCELL_X63_Y5_N0
\RegFile[18][6]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[18][6]~feeder_combout\ = ( \R.regWriteData\(6) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(6),
	combout => \RegFile[18][6]~feeder_combout\);

-- Location: FF_X63_Y5_N1
\RegFile[18][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][6]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][6]~q\);

-- Location: FF_X63_Y7_N37
\RegFile[19][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(6),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][6]~q\);

-- Location: LABCELL_X63_Y5_N45
\RegFile[16][6]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[16][6]~feeder_combout\ = \R.regWriteData\(6)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101010101010101010101010101010101010101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.regWriteData\(6),
	combout => \RegFile[16][6]~feeder_combout\);

-- Location: FF_X63_Y5_N46
\RegFile[16][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[16][6]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][6]~q\);

-- Location: MLABCELL_X65_Y8_N18
\Mux116~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux116~18_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[16][6]~q\))) # (\R.curInst\(20) & (\RegFile[17][6]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & (\RegFile[18][6]~q\)) # (\R.curInst\(20) & ((\RegFile[19][6]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[17][6]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[18][6]~q\,
	datad => \ALT_INV_RegFile[19][6]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][6]~q\,
	combout => \Mux116~18_combout\);

-- Location: FF_X68_Y7_N44
\RegFile[20][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(6),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][6]~q\);

-- Location: MLABCELL_X65_Y8_N36
\Mux116~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux116~5_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux116~18_combout\)))) # (\R.curInst\(22) & ((!\Mux116~18_combout\ & ((\RegFile[20][6]~q\))) # (\Mux116~18_combout\ & (\RegFile[21][6]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux116~18_combout\)))) # (\R.curInst\(22) & ((!\Mux116~18_combout\ & ((\RegFile[22][6]~q\))) # (\Mux116~18_combout\ & (\RegFile[23][6]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][6]~q\,
	datab => \ALT_INV_RegFile[23][6]~q\,
	datac => \ALT_INV_RegFile[22][6]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux116~18_combout\,
	datag => \ALT_INV_RegFile[20][6]~q\,
	combout => \Mux116~5_combout\);

-- Location: FF_X67_Y7_N2
\RegFile[3][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(6),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][6]~q\);

-- Location: FF_X68_Y7_N2
\RegFile[2][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(6),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][6]~q\);

-- Location: FF_X67_Y5_N40
\RegFile[4][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(6),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][6]~q\);

-- Location: FF_X63_Y7_N13
\RegFile[5][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(6),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][6]~q\);

-- Location: FF_X67_Y7_N25
\RegFile[7][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(6),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][6]~q\);

-- Location: FF_X67_Y7_N20
\RegFile[6][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(6),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][6]~q\);

-- Location: LABCELL_X67_Y7_N18
\Mux116~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux116~0_combout\ = ( \RegFile[6][6]~q\ & ( \R.curInst\(20) & ( (!\R.curInst\(21) & (\RegFile[5][6]~q\)) # (\R.curInst\(21) & ((\RegFile[7][6]~q\))) ) ) ) # ( !\RegFile[6][6]~q\ & ( \R.curInst\(20) & ( (!\R.curInst\(21) & (\RegFile[5][6]~q\)) # 
-- (\R.curInst\(21) & ((\RegFile[7][6]~q\))) ) ) ) # ( \RegFile[6][6]~q\ & ( !\R.curInst\(20) & ( (\R.curInst\(21)) # (\RegFile[4][6]~q\) ) ) ) # ( !\RegFile[6][6]~q\ & ( !\R.curInst\(20) & ( (\RegFile[4][6]~q\ & !\R.curInst\(21)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010100000000010101011111111100110011000011110011001100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[4][6]~q\,
	datab => \ALT_INV_RegFile[5][6]~q\,
	datac => \ALT_INV_RegFile[7][6]~q\,
	datad => \ALT_INV_R.curInst\(21),
	datae => \ALT_INV_RegFile[6][6]~q\,
	dataf => \ALT_INV_R.curInst\(20),
	combout => \Mux116~0_combout\);

-- Location: FF_X59_Y7_N50
\RegFile[1][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(6),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][6]~q\);

-- Location: LABCELL_X68_Y7_N0
\Mux116~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux116~26_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (\RegFile[1][6]~q\ & (\R.curInst\(20)))) # (\R.curInst\(22) & (((\Mux116~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (((\RegFile[2][6]~q\)))) # 
-- (\R.curInst\(20) & (\RegFile[3][6]~q\)))) # (\R.curInst\(22) & ((((\Mux116~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001100000011000100010000110011001111110011111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][6]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[2][6]~q\,
	datad => \ALT_INV_R.curInst\(20),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux116~0_combout\,
	datag => \ALT_INV_RegFile[1][6]~q\,
	combout => \Mux116~26_combout\);

-- Location: LABCELL_X64_Y6_N18
\RegFile[31][6]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[31][6]~feeder_combout\ = ( \R.regWriteData\(6) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(6),
	combout => \RegFile[31][6]~feeder_combout\);

-- Location: FF_X64_Y6_N19
\RegFile[31][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[31][6]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][6]~q\);

-- Location: MLABCELL_X52_Y7_N15
\RegFile[30][6]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[30][6]~feeder_combout\ = ( \R.regWriteData\(6) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(6),
	combout => \RegFile[30][6]~feeder_combout\);

-- Location: FF_X52_Y7_N16
\RegFile[30][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[30][6]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][6]~q\);

-- Location: FF_X59_Y7_N29
\RegFile[29][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(6),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][6]~q\);

-- Location: LABCELL_X64_Y6_N6
\RegFile[27][6]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[27][6]~feeder_combout\ = ( \R.regWriteData\(6) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(6),
	combout => \RegFile[27][6]~feeder_combout\);

-- Location: FF_X64_Y6_N8
\RegFile[27][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[27][6]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][6]~q\);

-- Location: FF_X59_Y7_N44
\RegFile[25][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(6),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][6]~q\);

-- Location: MLABCELL_X52_Y7_N39
\RegFile[26][6]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[26][6]~feeder_combout\ = ( \R.regWriteData\(6) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(6),
	combout => \RegFile[26][6]~feeder_combout\);

-- Location: FF_X52_Y7_N40
\RegFile[26][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[26][6]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][6]~q\);

-- Location: LABCELL_X64_Y6_N54
\RegFile[24][6]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[24][6]~feeder_combout\ = ( \R.regWriteData\(6) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(6),
	combout => \RegFile[24][6]~feeder_combout\);

-- Location: FF_X64_Y6_N56
\RegFile[24][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[24][6]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][6]~q\);

-- Location: MLABCELL_X59_Y7_N42
\Mux116~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux116~22_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[24][6]~q\))) # (\R.curInst\(20) & (\RegFile[25][6]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[26][6]~q\))) # (\R.curInst\(20) & (\RegFile[27][6]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[27][6]~q\,
	datab => \ALT_INV_RegFile[25][6]~q\,
	datac => \ALT_INV_RegFile[26][6]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][6]~q\,
	combout => \Mux116~22_combout\);

-- Location: FF_X65_Y9_N49
\RegFile[28][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(6),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][6]~q\);

-- Location: MLABCELL_X59_Y7_N27
\Mux116~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux116~9_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux116~22_combout\)))) # (\R.curInst\(22) & ((!\Mux116~22_combout\ & (\RegFile[28][6]~q\)) # (\Mux116~22_combout\ & ((\RegFile[29][6]~q\)))))) ) ) # ( \R.curInst\(21) & ( 
-- (!\R.curInst\(22) & ((((\Mux116~22_combout\))))) # (\R.curInst\(22) & (((!\Mux116~22_combout\ & ((\RegFile[30][6]~q\))) # (\Mux116~22_combout\ & (\RegFile[31][6]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111001100111111111101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][6]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[30][6]~q\,
	datad => \ALT_INV_RegFile[29][6]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux116~22_combout\,
	datag => \ALT_INV_RegFile[28][6]~q\,
	combout => \Mux116~9_combout\);

-- Location: FF_X64_Y7_N2
\RegFile[13][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(6),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][6]~q\);

-- Location: FF_X66_Y7_N26
\RegFile[15][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(6),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][6]~q\);

-- Location: FF_X61_Y7_N14
\RegFile[14][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(6),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][6]~q\);

-- Location: FF_X65_Y3_N14
\RegFile[9][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(6),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][6]~q\);

-- Location: MLABCELL_X65_Y3_N51
\RegFile[10][6]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[10][6]~feeder_combout\ = ( \R.regWriteData\(6) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(6),
	combout => \RegFile[10][6]~feeder_combout\);

-- Location: FF_X65_Y3_N53
\RegFile[10][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[10][6]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][6]~q\);

-- Location: FF_X65_Y3_N32
\RegFile[11][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(6),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][6]~q\);

-- Location: FF_X66_Y5_N44
\RegFile[8][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(6),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][6]~q\);

-- Location: MLABCELL_X65_Y3_N12
\Mux116~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux116~14_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[8][6]~q\))) # (\R.curInst\(20) & (\RegFile[9][6]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & (\RegFile[10][6]~q\)) # (\R.curInst\(20) & ((\RegFile[11][6]~q\)))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001110111011101110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[9][6]~q\,
	datac => \ALT_INV_RegFile[10][6]~q\,
	datad => \ALT_INV_RegFile[11][6]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][6]~q\,
	combout => \Mux116~14_combout\);

-- Location: LABCELL_X66_Y7_N39
\RegFile[12][6]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[12][6]~feeder_combout\ = ( \R.regWriteData\(6) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(6),
	combout => \RegFile[12][6]~feeder_combout\);

-- Location: FF_X66_Y7_N40
\RegFile[12][6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[12][6]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][6]~q\);

-- Location: LABCELL_X64_Y7_N0
\Mux116~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux116~1_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux116~14_combout\)))) # (\R.curInst\(22) & ((!\Mux116~14_combout\ & ((\RegFile[12][6]~q\))) # (\Mux116~14_combout\ & (\RegFile[13][6]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux116~14_combout\)))) # (\R.curInst\(22) & ((!\Mux116~14_combout\ & ((\RegFile[14][6]~q\))) # (\Mux116~14_combout\ & (\RegFile[15][6]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][6]~q\,
	datab => \ALT_INV_RegFile[15][6]~q\,
	datac => \ALT_INV_RegFile[14][6]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux116~14_combout\,
	datag => \ALT_INV_RegFile[12][6]~q\,
	combout => \Mux116~1_combout\);

-- Location: LABCELL_X74_Y7_N12
\Mux116~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux116~13_combout\ = ( \Mux116~9_combout\ & ( \Mux116~1_combout\ & ( ((!\R.curInst\(24) & ((\Mux116~26_combout\))) # (\R.curInst\(24) & (\Mux116~5_combout\))) # (\R.curInst\(23)) ) ) ) # ( !\Mux116~9_combout\ & ( \Mux116~1_combout\ & ( (!\R.curInst\(24) 
-- & (((\Mux116~26_combout\)) # (\R.curInst\(23)))) # (\R.curInst\(24) & (!\R.curInst\(23) & (\Mux116~5_combout\))) ) ) ) # ( \Mux116~9_combout\ & ( !\Mux116~1_combout\ & ( (!\R.curInst\(24) & (!\R.curInst\(23) & ((\Mux116~26_combout\)))) # (\R.curInst\(24) 
-- & (((\Mux116~5_combout\)) # (\R.curInst\(23)))) ) ) ) # ( !\Mux116~9_combout\ & ( !\Mux116~1_combout\ & ( (!\R.curInst\(23) & ((!\R.curInst\(24) & ((\Mux116~26_combout\))) # (\R.curInst\(24) & (\Mux116~5_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010010001100000101011001110100100110101011100011011110111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(24),
	datab => \ALT_INV_R.curInst\(23),
	datac => \ALT_INV_Mux116~5_combout\,
	datad => \ALT_INV_Mux116~26_combout\,
	datae => \ALT_INV_Mux116~9_combout\,
	dataf => \ALT_INV_Mux116~1_combout\,
	combout => \Mux116~13_combout\);

-- Location: LABCELL_X74_Y7_N45
\NxR.aluData2[6]~15\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[6]~15_combout\ = ( \Mux116~13_combout\ & ( (!\vAluSrc2~1_combout\) # ((\Equal4~1_combout\ & \Mux148~0_combout\)) ) ) # ( !\Mux116~13_combout\ & ( (\Equal4~1_combout\ & (\vAluSrc2~1_combout\ & \Mux148~0_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000101000000000000010111110000111101011111000011110101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Equal4~1_combout\,
	datac => \ALT_INV_vAluSrc2~1_combout\,
	datad => \ALT_INV_Mux148~0_combout\,
	dataf => \ALT_INV_Mux116~13_combout\,
	combout => \NxR.aluData2[6]~15_combout\);

-- Location: FF_X74_Y7_N56
\Add2~25_OTERM723_NEW_REG834\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \NxR.aluData2[6]~15_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Add2~25_OTERM723_OTERM835\);

-- Location: MLABCELL_X78_Y6_N21
\Add1~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~29_sumout\ = SUM(( \Add2~25_OTERM723_OTERM831\ ) + ( \Add2~25_OTERM723_OTERM829\ ) + ( \Add1~26\ ))
-- \Add1~30\ = CARRY(( \Add2~25_OTERM723_OTERM831\ ) + ( \Add2~25_OTERM723_OTERM829\ ) + ( \Add1~26\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add2~25_OTERM723_OTERM831\,
	datac => \ALT_INV_Add2~25_OTERM723_OTERM829\,
	cin => \Add1~26\,
	sumout => \Add1~29_sumout\,
	cout => \Add1~30\);

-- Location: MLABCELL_X78_Y6_N24
\Add1~33\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~33_sumout\ = SUM(( \Add2~33_OTERM719_OTERM827\ ) + ( \Add2~33_OTERM719_OTERM825\ ) + ( \Add1~30\ ))
-- \Add1~34\ = CARRY(( \Add2~33_OTERM719_OTERM827\ ) + ( \Add2~33_OTERM719_OTERM825\ ) + ( \Add1~30\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add2~33_OTERM719_OTERM825\,
	datad => \ALT_INV_Add2~33_OTERM719_OTERM827\,
	cin => \Add1~30\,
	sumout => \Add1~33_sumout\,
	cout => \Add1~34\);

-- Location: MLABCELL_X78_Y6_N27
\Add1~37\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~37_sumout\ = SUM(( \Add2~33_OTERM719_OTERM821\ ) + ( \Add2~33_OTERM719_OTERM823\ ) + ( \Add1~34\ ))
-- \Add1~38\ = CARRY(( \Add2~33_OTERM719_OTERM821\ ) + ( \Add2~33_OTERM719_OTERM823\ ) + ( \Add1~34\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Add2~33_OTERM719_OTERM823\,
	datad => \ALT_INV_Add2~33_OTERM719_OTERM821\,
	cin => \Add1~34\,
	sumout => \Add1~37_sumout\,
	cout => \Add1~38\);

-- Location: LABCELL_X80_Y3_N0
\Comb:vRegWriteData[9]~1_RESYN1080\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[9]~1_RESYN1080_BDD1081\ = ( \R.aluCalc~q\ & ( ((\R.aluOp.ALUOpSub~q\ & \Add2~37_sumout\)) # (\R.memToReg~q\) ) ) # ( !\R.aluCalc~q\ & ( (\R.memToReg~q\) # (\R.aluRes\(9)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011111100111111001111110011111100001111010111110000111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datab => \ALT_INV_R.aluRes\(9),
	datac => \ALT_INV_R.memToReg~q\,
	datad => \ALT_INV_Add2~37_sumout\,
	dataf => \ALT_INV_R.aluCalc~q\,
	combout => \Comb:vRegWriteData[9]~1_RESYN1080_BDD1081\);

-- Location: IOIBUF_X32_Y0_N18
\avm_d_readdata[17]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(17),
	o => \avm_d_readdata[17]~input_o\);

-- Location: LABCELL_X79_Y2_N48
\Comb:vRegWriteData[9]~1_RESYN1078\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[9]~1_RESYN1078_BDD1079\ = ( \avm_d_readdata[31]~input_o\ & ( \avm_d_readdata[17]~input_o\ & ( (!\R.memToReg~q\) # ((!\R.curInst\(12) & ((!\R.curInst\(14)))) # (\R.curInst\(12) & (!\R.curInst\(13)))) ) ) ) # ( 
-- !\avm_d_readdata[31]~input_o\ & ( \avm_d_readdata[17]~input_o\ & ( (!\R.memToReg~q\) # ((!\R.curInst\(13) & ((\R.curInst\(12)))) # (\R.curInst\(13) & (!\R.curInst\(14) & !\R.curInst\(12)))) ) ) ) # ( \avm_d_readdata[31]~input_o\ & ( 
-- !\avm_d_readdata[17]~input_o\ & ( (!\R.memToReg~q\) # ((!\R.curInst\(13) & (!\R.curInst\(14) & !\R.curInst\(12)))) ) ) ) # ( !\avm_d_readdata[31]~input_o\ & ( !\avm_d_readdata[17]~input_o\ & ( !\R.memToReg~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111100000000111111111000000011111111010010101111111111001010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(13),
	datab => \ALT_INV_R.curInst\(14),
	datac => \ALT_INV_R.curInst\(12),
	datad => \ALT_INV_R.memToReg~q\,
	datae => \ALT_INV_avm_d_readdata[31]~input_o\,
	dataf => \ALT_INV_avm_d_readdata[17]~input_o\,
	combout => \Comb:vRegWriteData[9]~1_RESYN1078_BDD1079\);

-- Location: LABCELL_X80_Y3_N36
\Comb:vRegWriteData[9]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[9]~1_combout\ = ( \Comb:vRegWriteData[9]~1_RESYN1080_BDD1081\ & ( \Comb:vRegWriteData[9]~1_RESYN1078_BDD1079\ ) ) # ( !\Comb:vRegWriteData[9]~1_RESYN1080_BDD1081\ & ( \Comb:vRegWriteData[9]~1_RESYN1078_BDD1079\ & ( (\R.aluCalc~q\ & 
-- ((!\Selector23~5_combout\) # ((\Add1~37_sumout\ & \R.aluOp.ALUOpAdd~q\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000001111000000011111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add1~37_sumout\,
	datab => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datac => \ALT_INV_R.aluCalc~q\,
	datad => \ALT_INV_Selector23~5_combout\,
	datae => \ALT_INV_Comb:vRegWriteData[9]~1_RESYN1080_BDD1081\,
	dataf => \ALT_INV_Comb:vRegWriteData[9]~1_RESYN1078_BDD1079\,
	combout => \Comb:vRegWriteData[9]~1_combout\);

-- Location: FF_X80_Y3_N5
\R.regWriteData[9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \R.regWriteData[9]~feeder_combout\,
	asdata => \Comb:vRegWriteData[9]~1_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(9));

-- Location: FF_X65_Y5_N14
\RegFile[13][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(9),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][9]~q\);

-- Location: FF_X65_Y5_N20
\RegFile[14][9]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(9),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][9]~DUPLICATE_q\);

-- Location: LABCELL_X64_Y3_N12
\Mux113~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux113~14_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & (\RegFile[8][9]~q\)) # (\R.curInst\(20) & ((\RegFile[9][9]~q\)))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & ((\RegFile[10][9]~q\))) # (\R.curInst\(20) & (\RegFile[11][9]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001010101111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[11][9]~q\,
	datac => \ALT_INV_RegFile[10][9]~q\,
	datad => \ALT_INV_RegFile[9][9]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][9]~q\,
	combout => \Mux113~14_combout\);

-- Location: MLABCELL_X65_Y5_N12
\Mux113~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux113~1_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux113~14_combout\))))) # (\R.curInst\(22) & (((!\Mux113~14_combout\ & ((\RegFile[12][9]~q\))) # (\Mux113~14_combout\ & (\RegFile[13][9]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux113~14_combout\)))) # (\R.curInst\(22) & ((!\Mux113~14_combout\ & (\RegFile[14][9]~DUPLICATE_q\)) # (\Mux113~14_combout\ & ((\RegFile[15][9]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][9]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[14][9]~DUPLICATE_q\,
	datad => \ALT_INV_RegFile[15][9]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux113~14_combout\,
	datag => \ALT_INV_RegFile[12][9]~q\,
	combout => \Mux113~1_combout\);

-- Location: LABCELL_X67_Y1_N12
\Mux113~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux113~22_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[24][9]~q\))) # (\R.curInst\(20) & (\RegFile[25][9]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & (\RegFile[26][9]~q\)) # (\R.curInst\(20) & ((\RegFile[27][9]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[25][9]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[26][9]~q\,
	datad => \ALT_INV_RegFile[27][9]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][9]~q\,
	combout => \Mux113~22_combout\);

-- Location: LABCELL_X64_Y1_N36
\Mux113~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux113~9_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux113~22_combout\))))) # (\R.curInst\(22) & (((!\Mux113~22_combout\ & ((\RegFile[28][9]~q\))) # (\Mux113~22_combout\ & (\RegFile[29][9]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux113~22_combout\)))) # (\R.curInst\(22) & ((!\Mux113~22_combout\ & (\RegFile[30][9]~q\)) # (\Mux113~22_combout\ & ((\RegFile[31][9]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[29][9]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[30][9]~q\,
	datad => \ALT_INV_RegFile[31][9]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux113~22_combout\,
	datag => \ALT_INV_RegFile[28][9]~q\,
	combout => \Mux113~9_combout\);

-- Location: LABCELL_X61_Y2_N42
\Mux113~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux113~0_combout\ = ( \RegFile[5][9]~q\ & ( \R.curInst\(21) & ( (!\R.curInst\(20) & (\RegFile[6][9]~q\)) # (\R.curInst\(20) & ((\RegFile[7][9]~q\))) ) ) ) # ( !\RegFile[5][9]~q\ & ( \R.curInst\(21) & ( (!\R.curInst\(20) & (\RegFile[6][9]~q\)) # 
-- (\R.curInst\(20) & ((\RegFile[7][9]~q\))) ) ) ) # ( \RegFile[5][9]~q\ & ( !\R.curInst\(21) & ( (\RegFile[4][9]~q\) # (\R.curInst\(20)) ) ) ) # ( !\RegFile[5][9]~q\ & ( !\R.curInst\(21) & ( (!\R.curInst\(20) & \RegFile[4][9]~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011110000000011111111111101010011010100110101001101010011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[6][9]~q\,
	datab => \ALT_INV_RegFile[7][9]~q\,
	datac => \ALT_INV_R.curInst\(20),
	datad => \ALT_INV_RegFile[4][9]~q\,
	datae => \ALT_INV_RegFile[5][9]~q\,
	dataf => \ALT_INV_R.curInst\(21),
	combout => \Mux113~0_combout\);

-- Location: LABCELL_X64_Y5_N12
\Mux113~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux113~26_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (\R.curInst\(20) & (\RegFile[1][9]~q\))) # (\R.curInst\(22) & (((\Mux113~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (((\RegFile[2][9]~q\)))) # 
-- (\R.curInst\(20) & (\RegFile[3][9]~q\)))) # (\R.curInst\(22) & ((((\Mux113~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000000000110110000000000000101111111110001101111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(20),
	datab => \ALT_INV_RegFile[3][9]~q\,
	datac => \ALT_INV_RegFile[2][9]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux113~0_combout\,
	datag => \ALT_INV_RegFile[1][9]~q\,
	combout => \Mux113~26_combout\);

-- Location: FF_X64_Y4_N1
\RegFile[22][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[22][9]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][9]~q\);

-- Location: FF_X57_Y5_N11
\RegFile[17][9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(9),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][9]~q\);

-- Location: LABCELL_X57_Y5_N48
\Mux113~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux113~18_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & (\RegFile[16][9]~q\)) # (\R.curInst\(20) & ((\RegFile[17][9]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & ((\RegFile[18][9]~q\))) # (\R.curInst\(20) & (\RegFile[19][9]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110000110011111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[19][9]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[18][9]~q\,
	datad => \ALT_INV_RegFile[17][9]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][9]~q\,
	combout => \Mux113~18_combout\);

-- Location: LABCELL_X64_Y5_N3
\Mux113~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux113~5_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux113~18_combout\)))) # (\R.curInst\(22) & ((!\Mux113~18_combout\ & (\RegFile[20][9]~q\)) # (\Mux113~18_combout\ & ((\RegFile[21][9]~q\)))))) ) ) # ( \R.curInst\(21) & ( 
-- (!\R.curInst\(22) & ((((\Mux113~18_combout\))))) # (\R.curInst\(22) & (((!\Mux113~18_combout\ & ((\RegFile[22][9]~q\))) # (\Mux113~18_combout\ & (\RegFile[23][9]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111001100111111111101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[23][9]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[22][9]~q\,
	datad => \ALT_INV_RegFile[21][9]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux113~18_combout\,
	datag => \ALT_INV_RegFile[20][9]~q\,
	combout => \Mux113~5_combout\);

-- Location: MLABCELL_X65_Y5_N21
\Mux113~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux113~13_combout\ = ( \Mux113~26_combout\ & ( \Mux113~5_combout\ & ( (!\R.curInst\(23)) # ((!\R.curInst\(24) & (\Mux113~1_combout\)) # (\R.curInst\(24) & ((\Mux113~9_combout\)))) ) ) ) # ( !\Mux113~26_combout\ & ( \Mux113~5_combout\ & ( 
-- (!\R.curInst\(23) & (((\R.curInst\(24))))) # (\R.curInst\(23) & ((!\R.curInst\(24) & (\Mux113~1_combout\)) # (\R.curInst\(24) & ((\Mux113~9_combout\))))) ) ) ) # ( \Mux113~26_combout\ & ( !\Mux113~5_combout\ & ( (!\R.curInst\(23) & (((!\R.curInst\(24))))) 
-- # (\R.curInst\(23) & ((!\R.curInst\(24) & (\Mux113~1_combout\)) # (\R.curInst\(24) & ((\Mux113~9_combout\))))) ) ) ) # ( !\Mux113~26_combout\ & ( !\Mux113~5_combout\ & ( (\R.curInst\(23) & ((!\R.curInst\(24) & (\Mux113~1_combout\)) # (\R.curInst\(24) & 
-- ((\Mux113~9_combout\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100000101101110110000010100010001101011111011101110101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(23),
	datab => \ALT_INV_Mux113~1_combout\,
	datac => \ALT_INV_Mux113~9_combout\,
	datad => \ALT_INV_R.curInst\(24),
	datae => \ALT_INV_Mux113~26_combout\,
	dataf => \ALT_INV_Mux113~5_combout\,
	combout => \Mux113~13_combout\);

-- Location: LABCELL_X74_Y7_N0
\NxR.aluData2[9]~12\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[9]~12_combout\ = ( \Mux113~13_combout\ & ( (!\vAluSrc2~1_combout\) # ((\Equal4~1_combout\ & \Mux145~0_combout\)) ) ) # ( !\Mux113~13_combout\ & ( (\vAluSrc2~1_combout\ & (\Equal4~1_combout\ & \Mux145~0_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000011000000000000001111001100110011111100110011001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_vAluSrc2~1_combout\,
	datac => \ALT_INV_Equal4~1_combout\,
	datad => \ALT_INV_Mux145~0_combout\,
	dataf => \ALT_INV_Mux113~13_combout\,
	combout => \NxR.aluData2[9]~12_combout\);

-- Location: FF_X74_Y7_N22
\Add2~33_OTERM719_NEW_REG822\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \NxR.aluData2[9]~12_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Add2~33_OTERM719_OTERM823\);

-- Location: MLABCELL_X78_Y6_N30
\Add1~41\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~41_sumout\ = SUM(( \Add2~41_OTERM715_OTERM817\ ) + ( \Add2~41_OTERM715_OTERM819\ ) + ( \Add1~38\ ))
-- \Add1~42\ = CARRY(( \Add2~41_OTERM715_OTERM817\ ) + ( \Add2~41_OTERM715_OTERM819\ ) + ( \Add1~38\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Add2~41_OTERM715_OTERM819\,
	datad => \ALT_INV_Add2~41_OTERM715_OTERM817\,
	cin => \Add1~38\,
	sumout => \Add1~41_sumout\,
	cout => \Add1~42\);

-- Location: MLABCELL_X78_Y6_N33
\Add1~45\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~45_sumout\ = SUM(( \R.aluData1\(11) ) + ( \R.aluData2\(11) ) + ( \Add1~42\ ))
-- \Add1~46\ = CARRY(( \R.aluData1\(11) ) + ( \R.aluData2\(11) ) + ( \Add1~42\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData1\(11),
	dataf => \ALT_INV_R.aluData2\(11),
	cin => \Add1~42\,
	sumout => \Add1~45_sumout\,
	cout => \Add1~46\);

-- Location: MLABCELL_X78_Y6_N39
\Add1~53\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~53_sumout\ = SUM(( \R.aluData1\(13) ) + ( \R.aluData2\(13) ) + ( \Add1~50\ ))
-- \Add1~54\ = CARRY(( \R.aluData1\(13) ) + ( \R.aluData2\(13) ) + ( \Add1~50\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(13),
	datad => \ALT_INV_R.aluData1\(13),
	cin => \Add1~50\,
	sumout => \Add1~53_sumout\,
	cout => \Add1~54\);

-- Location: IOIBUF_X60_Y0_N52
\avm_d_readdata[22]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(22),
	o => \avm_d_readdata[22]~input_o\);

-- Location: LABCELL_X79_Y2_N45
\Comb:vRegWriteData[14]~1_RESYN1094\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[14]~1_RESYN1094_BDD1095\ = ( \R.curInst\(13) & ( \R.curInst\(12) & ( !\R.memToReg~q\ ) ) ) # ( !\R.curInst\(13) & ( \R.curInst\(12) & ( (!\R.memToReg~q\) # (\avm_d_readdata[22]~input_o\) ) ) ) # ( \R.curInst\(13) & ( !\R.curInst\(12) & 
-- ( (!\R.memToReg~q\) # ((!\R.curInst\(14) & \avm_d_readdata[22]~input_o\)) ) ) ) # ( !\R.curInst\(13) & ( !\R.curInst\(12) & ( (!\R.memToReg~q\) # ((!\R.curInst\(14) & \avm_d_readdata[31]~input_o\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111001011110010111100001111101011110000111111111111000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(14),
	datab => \ALT_INV_avm_d_readdata[31]~input_o\,
	datac => \ALT_INV_R.memToReg~q\,
	datad => \ALT_INV_avm_d_readdata[22]~input_o\,
	datae => \ALT_INV_R.curInst\(13),
	dataf => \ALT_INV_R.curInst\(12),
	combout => \Comb:vRegWriteData[14]~1_RESYN1094_BDD1095\);

-- Location: LABCELL_X80_Y3_N30
\Comb:vRegWriteData[14]~1_RESYN1096\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[14]~1_RESYN1096_BDD1097\ = ( \R.aluCalc~q\ & ( ((\R.aluOp.ALUOpSub~q\ & \Add2~57_sumout\)) # (\R.memToReg~q\) ) ) # ( !\R.aluCalc~q\ & ( (\R.aluRes\(14)) # (\R.memToReg~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0111011101110111011101110111011101010101010111110101010101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.memToReg~q\,
	datab => \ALT_INV_R.aluRes\(14),
	datac => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datad => \ALT_INV_Add2~57_sumout\,
	dataf => \ALT_INV_R.aluCalc~q\,
	combout => \Comb:vRegWriteData[14]~1_RESYN1096_BDD1097\);

-- Location: LABCELL_X80_Y3_N54
\Comb:vRegWriteData[14]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[14]~1_combout\ = ( \Comb:vRegWriteData[14]~1_RESYN1094_BDD1095\ & ( \Comb:vRegWriteData[14]~1_RESYN1096_BDD1097\ ) ) # ( \Comb:vRegWriteData[14]~1_RESYN1094_BDD1095\ & ( !\Comb:vRegWriteData[14]~1_RESYN1096_BDD1097\ & ( (\R.aluCalc~q\ 
-- & ((!\Selector18~3_combout\) # ((\Add1~57_sumout\ & \R.aluOp.ALUOpAdd~q\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000001100000011000100000000000000001111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add1~57_sumout\,
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_Selector18~3_combout\,
	datad => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datae => \ALT_INV_Comb:vRegWriteData[14]~1_RESYN1094_BDD1095\,
	dataf => \ALT_INV_Comb:vRegWriteData[14]~1_RESYN1096_BDD1097\,
	combout => \Comb:vRegWriteData[14]~1_combout\);

-- Location: FF_X80_Y3_N35
\R.regWriteData[14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \R.regWriteData[14]~feeder_combout\,
	asdata => \Comb:vRegWriteData[14]~1_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(14));

-- Location: FF_X66_Y6_N2
\RegFile[29][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(14),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][14]~q\);

-- Location: LABCELL_X57_Y6_N33
\RegFile[30][14]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[30][14]~feeder_combout\ = ( \R.regWriteData\(14) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(14),
	combout => \RegFile[30][14]~feeder_combout\);

-- Location: FF_X57_Y6_N34
\RegFile[30][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[30][14]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][14]~q\);

-- Location: FF_X64_Y6_N2
\RegFile[31][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(14),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][14]~q\);

-- Location: FF_X66_Y6_N20
\RegFile[25][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(14),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][14]~q\);

-- Location: LABCELL_X64_Y6_N36
\RegFile[27][14]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[27][14]~feeder_combout\ = ( \R.regWriteData\(14) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(14),
	combout => \RegFile[27][14]~feeder_combout\);

-- Location: FF_X64_Y6_N37
\RegFile[27][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[27][14]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][14]~q\);

-- Location: LABCELL_X57_Y6_N36
\RegFile[26][14]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[26][14]~feeder_combout\ = ( \R.regWriteData\(14) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(14),
	combout => \RegFile[26][14]~feeder_combout\);

-- Location: FF_X57_Y6_N37
\RegFile[26][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[26][14]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][14]~q\);

-- Location: LABCELL_X64_Y6_N45
\RegFile[24][14]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[24][14]~feeder_combout\ = ( \R.regWriteData\(14) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(14),
	combout => \RegFile[24][14]~feeder_combout\);

-- Location: FF_X64_Y6_N46
\RegFile[24][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[24][14]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][14]~q\);

-- Location: LABCELL_X66_Y6_N18
\Mux108~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux108~22_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[24][14]~q\))) # (\R.curInst\(20) & (\RegFile[25][14]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[26][14]~q\))) # (\R.curInst\(20) & (\RegFile[27][14]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[25][14]~q\,
	datab => \ALT_INV_RegFile[27][14]~q\,
	datac => \ALT_INV_RegFile[26][14]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][14]~q\,
	combout => \Mux108~22_combout\);

-- Location: FF_X65_Y9_N22
\RegFile[28][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(14),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][14]~q\);

-- Location: LABCELL_X66_Y6_N0
\Mux108~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux108~9_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux108~22_combout\))))) # (\R.curInst\(22) & (((!\Mux108~22_combout\ & ((\RegFile[28][14]~q\))) # (\Mux108~22_combout\ & (\RegFile[29][14]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux108~22_combout\)))) # (\R.curInst\(22) & ((!\Mux108~22_combout\ & (\RegFile[30][14]~q\)) # (\Mux108~22_combout\ & ((\RegFile[31][14]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[29][14]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[30][14]~q\,
	datad => \ALT_INV_RegFile[31][14]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux108~22_combout\,
	datag => \ALT_INV_RegFile[28][14]~q\,
	combout => \Mux108~9_combout\);

-- Location: LABCELL_X68_Y6_N54
\RegFile[21][14]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[21][14]~feeder_combout\ = ( \R.regWriteData\(14) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(14),
	combout => \RegFile[21][14]~feeder_combout\);

-- Location: FF_X68_Y6_N56
\RegFile[21][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[21][14]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][14]~q\);

-- Location: FF_X64_Y4_N59
\RegFile[22][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(14),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][14]~q\);

-- Location: FF_X64_Y2_N38
\RegFile[23][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(14),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][14]~q\);

-- Location: FF_X65_Y2_N38
\RegFile[17][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(14),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][14]~q\);

-- Location: FF_X64_Y2_N44
\RegFile[19][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(14),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][14]~q\);

-- Location: FF_X57_Y2_N7
\RegFile[18][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(14),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][14]~q\);

-- Location: FF_X57_Y2_N40
\RegFile[16][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(14),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][14]~q\);

-- Location: MLABCELL_X65_Y2_N36
\Mux108~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux108~18_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[16][14]~q\))) # (\R.curInst\(20) & (\RegFile[17][14]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[18][14]~q\))) # (\R.curInst\(20) & (\RegFile[19][14]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[17][14]~q\,
	datab => \ALT_INV_RegFile[19][14]~q\,
	datac => \ALT_INV_RegFile[18][14]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][14]~q\,
	combout => \Mux108~18_combout\);

-- Location: LABCELL_X68_Y6_N24
\RegFile[20][14]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[20][14]~feeder_combout\ = ( \R.regWriteData\(14) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(14),
	combout => \RegFile[20][14]~feeder_combout\);

-- Location: FF_X68_Y6_N25
\RegFile[20][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[20][14]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][14]~q\);

-- Location: LABCELL_X68_Y6_N48
\Mux108~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux108~5_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux108~18_combout\))))) # (\R.curInst\(22) & (((!\Mux108~18_combout\ & ((\RegFile[20][14]~q\))) # (\Mux108~18_combout\ & (\RegFile[21][14]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux108~18_combout\)))) # (\R.curInst\(22) & ((!\Mux108~18_combout\ & (\RegFile[22][14]~q\)) # (\Mux108~18_combout\ & ((\RegFile[23][14]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][14]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[22][14]~q\,
	datad => \ALT_INV_RegFile[23][14]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux108~18_combout\,
	datag => \ALT_INV_RegFile[20][14]~q\,
	combout => \Mux108~5_combout\);

-- Location: FF_X62_Y8_N32
\RegFile[3][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(14),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][14]~q\);

-- Location: FF_X61_Y4_N56
\RegFile[2][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(14),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][14]~q\);

-- Location: FF_X62_Y8_N14
\RegFile[7][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(14),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][14]~q\);

-- Location: LABCELL_X62_Y8_N54
\RegFile[5][14]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[5][14]~feeder_combout\ = ( \R.regWriteData\(14) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(14),
	combout => \RegFile[5][14]~feeder_combout\);

-- Location: FF_X62_Y8_N55
\RegFile[5][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[5][14]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][14]~q\);

-- Location: LABCELL_X56_Y4_N45
\RegFile[4][14]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[4][14]~feeder_combout\ = ( \R.regWriteData\(14) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(14),
	combout => \RegFile[4][14]~feeder_combout\);

-- Location: FF_X56_Y4_N46
\RegFile[4][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[4][14]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][14]~q\);

-- Location: FF_X61_Y4_N19
\RegFile[6][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(14),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][14]~q\);

-- Location: LABCELL_X61_Y4_N18
\Mux108~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux108~0_combout\ = ( \RegFile[6][14]~q\ & ( \R.curInst\(20) & ( (!\R.curInst\(21) & ((\RegFile[5][14]~q\))) # (\R.curInst\(21) & (\RegFile[7][14]~q\)) ) ) ) # ( !\RegFile[6][14]~q\ & ( \R.curInst\(20) & ( (!\R.curInst\(21) & ((\RegFile[5][14]~q\))) # 
-- (\R.curInst\(21) & (\RegFile[7][14]~q\)) ) ) ) # ( \RegFile[6][14]~q\ & ( !\R.curInst\(20) & ( (\R.curInst\(21)) # (\RegFile[4][14]~q\) ) ) ) # ( !\RegFile[6][14]~q\ & ( !\R.curInst\(20) & ( (\RegFile[4][14]~q\ & !\R.curInst\(21)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100000000000011111111111100110011010101010011001101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[7][14]~q\,
	datab => \ALT_INV_RegFile[5][14]~q\,
	datac => \ALT_INV_RegFile[4][14]~q\,
	datad => \ALT_INV_R.curInst\(21),
	datae => \ALT_INV_RegFile[6][14]~q\,
	dataf => \ALT_INV_R.curInst\(20),
	combout => \Mux108~0_combout\);

-- Location: MLABCELL_X59_Y7_N57
\RegFile[1][14]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[1][14]~feeder_combout\ = ( \R.regWriteData\(14) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(14),
	combout => \RegFile[1][14]~feeder_combout\);

-- Location: FF_X59_Y7_N59
\RegFile[1][14]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[1][14]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][14]~DUPLICATE_q\);

-- Location: LABCELL_X61_Y4_N54
\Mux108~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux108~26_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (\R.curInst\(20) & (\RegFile[1][14]~DUPLICATE_q\))) # (\R.curInst\(22) & (((\Mux108~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & 
-- (((\RegFile[2][14]~q\)))) # (\R.curInst\(20) & (\RegFile[3][14]~q\)))) # (\R.curInst\(22) & ((((\Mux108~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000000000110110000000000000101111111110001101111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(20),
	datab => \ALT_INV_RegFile[3][14]~q\,
	datac => \ALT_INV_RegFile[2][14]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux108~0_combout\,
	datag => \ALT_INV_RegFile[1][14]~DUPLICATE_q\,
	combout => \Mux108~26_combout\);

-- Location: FF_X63_Y6_N50
\RegFile[15][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(14),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][14]~q\);

-- Location: FF_X67_Y8_N26
\RegFile[13][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(14),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][14]~q\);

-- Location: LABCELL_X67_Y8_N12
\RegFile[14][14]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[14][14]~feeder_combout\ = ( \R.regWriteData\(14) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(14),
	combout => \RegFile[14][14]~feeder_combout\);

-- Location: FF_X67_Y8_N13
\RegFile[14][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[14][14]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][14]~q\);

-- Location: FF_X67_Y8_N44
\RegFile[9][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(14),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][14]~q\);

-- Location: LABCELL_X64_Y8_N15
\RegFile[10][14]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[10][14]~feeder_combout\ = ( \R.regWriteData\(14) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(14),
	combout => \RegFile[10][14]~feeder_combout\);

-- Location: FF_X64_Y8_N16
\RegFile[10][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[10][14]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][14]~q\);

-- Location: FF_X63_Y6_N32
\RegFile[11][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(14),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][14]~q\);

-- Location: LABCELL_X63_Y6_N54
\RegFile[8][14]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[8][14]~feeder_combout\ = ( \R.regWriteData\(14) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(14),
	combout => \RegFile[8][14]~feeder_combout\);

-- Location: FF_X63_Y6_N56
\RegFile[8][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[8][14]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][14]~q\);

-- Location: LABCELL_X67_Y8_N42
\Mux108~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux108~14_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[8][14]~q\))) # (\R.curInst\(20) & (\RegFile[9][14]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & (\RegFile[10][14]~q\)) # (\R.curInst\(20) & ((\RegFile[11][14]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][14]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[10][14]~q\,
	datad => \ALT_INV_RegFile[11][14]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][14]~q\,
	combout => \Mux108~14_combout\);

-- Location: LABCELL_X66_Y7_N3
\RegFile[12][14]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[12][14]~feeder_combout\ = ( \R.regWriteData\(14) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(14),
	combout => \RegFile[12][14]~feeder_combout\);

-- Location: FF_X66_Y7_N4
\RegFile[12][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[12][14]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][14]~q\);

-- Location: LABCELL_X67_Y8_N24
\Mux108~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux108~1_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux108~14_combout\)))) # (\R.curInst\(22) & ((!\Mux108~14_combout\ & ((\RegFile[12][14]~q\))) # (\Mux108~14_combout\ & (\RegFile[13][14]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux108~14_combout\)))) # (\R.curInst\(22) & ((!\Mux108~14_combout\ & ((\RegFile[14][14]~q\))) # (\Mux108~14_combout\ & (\RegFile[15][14]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][14]~q\,
	datab => \ALT_INV_RegFile[13][14]~q\,
	datac => \ALT_INV_RegFile[14][14]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux108~14_combout\,
	datag => \ALT_INV_RegFile[12][14]~q\,
	combout => \Mux108~1_combout\);

-- Location: LABCELL_X75_Y6_N48
\Mux108~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux108~13_combout\ = ( \Mux108~26_combout\ & ( \Mux108~1_combout\ & ( (!\R.curInst\(24)) # ((!\R.curInst\(23) & ((\Mux108~5_combout\))) # (\R.curInst\(23) & (\Mux108~9_combout\))) ) ) ) # ( !\Mux108~26_combout\ & ( \Mux108~1_combout\ & ( 
-- (!\R.curInst\(23) & (\R.curInst\(24) & ((\Mux108~5_combout\)))) # (\R.curInst\(23) & ((!\R.curInst\(24)) # ((\Mux108~9_combout\)))) ) ) ) # ( \Mux108~26_combout\ & ( !\Mux108~1_combout\ & ( (!\R.curInst\(23) & ((!\R.curInst\(24)) # 
-- ((\Mux108~5_combout\)))) # (\R.curInst\(23) & (\R.curInst\(24) & (\Mux108~9_combout\))) ) ) ) # ( !\Mux108~26_combout\ & ( !\Mux108~1_combout\ & ( (\R.curInst\(24) & ((!\R.curInst\(23) & ((\Mux108~5_combout\))) # (\R.curInst\(23) & (\Mux108~9_combout\)))) 
-- ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000100100011100010011010101101000101011001111100110111101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(23),
	datab => \ALT_INV_R.curInst\(24),
	datac => \ALT_INV_Mux108~9_combout\,
	datad => \ALT_INV_Mux108~5_combout\,
	datae => \ALT_INV_Mux108~26_combout\,
	dataf => \ALT_INV_Mux108~1_combout\,
	combout => \Mux108~13_combout\);

-- Location: LABCELL_X75_Y6_N33
\NxR.aluData2[14]~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[14]~7_combout\ = ( \Mux108~13_combout\ & ( (!\vAluSrc2~1_combout\) # ((\Mux140~0_combout\ & \Equal4~1_combout\)) ) ) # ( !\Mux108~13_combout\ & ( (\Mux140~0_combout\ & (\vAluSrc2~1_combout\ & \Equal4~1_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000101000000000000010111110000111101011111000011110101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux140~0_combout\,
	datac => \ALT_INV_vAluSrc2~1_combout\,
	datad => \ALT_INV_Equal4~1_combout\,
	dataf => \ALT_INV_Mux108~13_combout\,
	combout => \NxR.aluData2[14]~7_combout\);

-- Location: FF_X75_Y6_N10
\Add2~57_OTERM707_NEW_REG814\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \NxR.aluData2[14]~7_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Add2~57_OTERM707_OTERM815\);

-- Location: LABCELL_X77_Y7_N30
\ShiftRight1~54\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~54_combout\ = ( \ShiftRight1~32_OTERM21\ & ( \ShiftRight1~31_OTERM45\ & ( ((!\R.aluData2\(2) & (\ShiftRight1~37_OTERM283\)) # (\R.aluData2\(2) & ((\ShiftRight1~30_OTERM39\)))) # (\R.aluData2\(3)) ) ) ) # ( !\ShiftRight1~32_OTERM21\ & ( 
-- \ShiftRight1~31_OTERM45\ & ( (!\R.aluData2\(2) & (((\R.aluData2\(3))) # (\ShiftRight1~37_OTERM283\))) # (\R.aluData2\(2) & (((\ShiftRight1~30_OTERM39\ & !\R.aluData2\(3))))) ) ) ) # ( \ShiftRight1~32_OTERM21\ & ( !\ShiftRight1~31_OTERM45\ & ( 
-- (!\R.aluData2\(2) & (\ShiftRight1~37_OTERM283\ & ((!\R.aluData2\(3))))) # (\R.aluData2\(2) & (((\R.aluData2\(3)) # (\ShiftRight1~30_OTERM39\)))) ) ) ) # ( !\ShiftRight1~32_OTERM21\ & ( !\ShiftRight1~31_OTERM45\ & ( (!\R.aluData2\(3) & ((!\R.aluData2\(2) & 
-- (\ShiftRight1~37_OTERM283\)) # (\R.aluData2\(2) & ((\ShiftRight1~30_OTERM39\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100011100000000010001110011001101000111110011000100011111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~37_OTERM283\,
	datab => \ALT_INV_R.aluData2\(2),
	datac => \ALT_INV_ShiftRight1~30_OTERM39\,
	datad => \ALT_INV_R.aluData2\(3),
	datae => \ALT_INV_ShiftRight1~32_OTERM21\,
	dataf => \ALT_INV_ShiftRight1~31_OTERM45\,
	combout => \ShiftRight1~54_combout\);

-- Location: LABCELL_X77_Y7_N24
\Selector17~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector17~1_combout\ = ( \R.aluData1\(15) & ( \R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( (!\R.aluOp.ALUOpXor~DUPLICATE_q\ & (!\R.aluData2\(15) & !\R.aluOp.ALUOpOr~q\)) ) ) ) # ( !\R.aluData1\(15) & ( \R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( (!\R.aluData2\(15)) # 
-- ((!\R.aluOp.ALUOpXor~DUPLICATE_q\ & !\R.aluOp.ALUOpOr~q\)) ) ) ) # ( \R.aluData1\(15) & ( !\R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( (!\R.aluOp.ALUOpOr~q\ & ((!\R.aluOp.ALUOpXor~DUPLICATE_q\) # (\R.aluData2\(15)))) ) ) ) # ( !\R.aluData1\(15) & ( 
-- !\R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( (!\R.aluData2\(15)) # ((!\R.aluOp.ALUOpXor~DUPLICATE_q\ & !\R.aluOp.ALUOpOr~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1110110011101100101100001011000011101100111011001000000010000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpXor~DUPLICATE_q\,
	datab => \ALT_INV_R.aluData2\(15),
	datac => \ALT_INV_R.aluOp.ALUOpOr~q\,
	datae => \ALT_INV_R.aluData1\(15),
	dataf => \ALT_INV_R.aluOp.ALUOpAnd~DUPLICATE_q\,
	combout => \Selector17~1_combout\);

-- Location: LABCELL_X77_Y7_N18
\Selector17~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector17~2_combout\ = ( \Selector31~7_OTERM383\ & ( (\Selector17~1_combout\ & (!\Selector17~0_OTERM391\ & ((!\ShiftRight0~4_OTERM31\) # (\ShiftRight0~7_OTERM233DUPLICATE_q\)))) ) ) # ( !\Selector31~7_OTERM383\ & ( (\Selector17~1_combout\ & 
-- !\Selector17~0_OTERM391\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100000000000011110000000000001011000000000000101100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight0~4_OTERM31\,
	datab => \ALT_INV_ShiftRight0~7_OTERM233DUPLICATE_q\,
	datac => \ALT_INV_Selector17~1_combout\,
	datad => \ALT_INV_Selector17~0_OTERM391\,
	dataf => \ALT_INV_Selector31~7_OTERM383\,
	combout => \Selector17~2_combout\);

-- Location: LABCELL_X79_Y8_N24
\Selector17~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector17~3_combout\ = ( \R.aluOp.ALUOpSLL~q\ & ( \ShiftLeft0~23_combout\ & ( (!\R.aluData2\(4)) # (!\Selector17~2_combout\) ) ) ) # ( !\R.aluOp.ALUOpSLL~q\ & ( \ShiftLeft0~23_combout\ & ( (!\Selector17~2_combout\) # ((\ShiftRight1~54_combout\ & 
-- (\Selector31~0_OTERM349\ & !\R.aluData2\(4)))) ) ) ) # ( \R.aluOp.ALUOpSLL~q\ & ( !\ShiftLeft0~23_combout\ & ( (!\Selector17~2_combout\) # ((\ShiftRight1~54_combout\ & (\Selector31~0_OTERM349\ & !\R.aluData2\(4)))) ) ) ) # ( !\R.aluOp.ALUOpSLL~q\ & ( 
-- !\ShiftLeft0~23_combout\ & ( (!\Selector17~2_combout\) # ((\ShiftRight1~54_combout\ & (\Selector31~0_OTERM349\ & !\R.aluData2\(4)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111100010000111111110001000011111111000100001111111111110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~54_combout\,
	datab => \ALT_INV_Selector31~0_OTERM349\,
	datac => \ALT_INV_R.aluData2\(4),
	datad => \ALT_INV_Selector17~2_combout\,
	datae => \ALT_INV_R.aluOp.ALUOpSLL~q\,
	dataf => \ALT_INV_ShiftLeft0~23_combout\,
	combout => \Selector17~3_combout\);

-- Location: LABCELL_X80_Y6_N0
\Selector17~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector17~5_combout\ = ( \Selector17~3_combout\ ) # ( !\Selector17~3_combout\ & ( (!\Add2~61_sumout\ & (((\Add1~61_sumout\ & \R.aluOp.ALUOpAdd~q\)))) # (\Add2~61_sumout\ & (((\Add1~61_sumout\ & \R.aluOp.ALUOpAdd~q\)) # (\R.aluOp.ALUOpSub~q\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100011111000100010001111111111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add2~61_sumout\,
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_Add1~61_sumout\,
	datad => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	dataf => \ALT_INV_Selector17~3_combout\,
	combout => \Selector17~5_combout\);

-- Location: FF_X80_Y6_N2
\R.aluRes[15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector17~5_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(15));

-- Location: LABCELL_X80_Y6_N3
\Comb:vRegWriteData[15]~1_RESYN1048\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[15]~1_RESYN1048_BDD1049\ = ( \R.memToReg~q\ ) # ( !\R.memToReg~q\ & ( (!\R.aluCalc~q\ & (((\R.aluRes\(15))))) # (\R.aluCalc~q\ & (\Add2~61_sumout\ & (\R.aluOp.ALUOpSub~q\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000111110001000000011111000111111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add2~61_sumout\,
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_R.aluCalc~q\,
	datad => \ALT_INV_R.aluRes\(15),
	dataf => \ALT_INV_R.memToReg~q\,
	combout => \Comb:vRegWriteData[15]~1_RESYN1048_BDD1049\);

-- Location: LABCELL_X80_Y2_N15
\Comb:vRegWriteData[15]~1_RESYN1046\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[15]~1_RESYN1046_BDD1047\ = ( \R.curInst\(13) & ( \R.curInst\(12) & ( !\R.memToReg~q\ ) ) ) # ( !\R.curInst\(13) & ( \R.curInst\(12) & ( (!\R.memToReg~q\) # (\avm_d_readdata[23]~input_o\) ) ) ) # ( \R.curInst\(13) & ( !\R.curInst\(12) & 
-- ( (!\R.memToReg~q\) # ((\avm_d_readdata[23]~input_o\ & !\R.curInst\(14))) ) ) ) # ( !\R.curInst\(13) & ( !\R.curInst\(12) & ( (!\R.memToReg~q\) # ((\avm_d_readdata[31]~input_o\ & !\R.curInst\(14))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111101010000111111110011000011111111001100111111111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_avm_d_readdata[31]~input_o\,
	datab => \ALT_INV_avm_d_readdata[23]~input_o\,
	datac => \ALT_INV_R.curInst\(14),
	datad => \ALT_INV_R.memToReg~q\,
	datae => \ALT_INV_R.curInst\(13),
	dataf => \ALT_INV_R.curInst\(12),
	combout => \Comb:vRegWriteData[15]~1_RESYN1046_BDD1047\);

-- Location: LABCELL_X80_Y6_N48
\Comb:vRegWriteData[15]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[15]~1_combout\ = ( \R.aluCalc~q\ & ( \Comb:vRegWriteData[15]~1_RESYN1046_BDD1047\ & ( (((\R.aluOp.ALUOpAdd~q\ & \Add1~61_sumout\)) # (\Selector17~3_combout\)) # (\Comb:vRegWriteData[15]~1_RESYN1048_BDD1049\) ) ) ) # ( !\R.aluCalc~q\ & 
-- ( \Comb:vRegWriteData[15]~1_RESYN1046_BDD1047\ & ( \Comb:vRegWriteData[15]~1_RESYN1048_BDD1049\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000001010101010101010101011111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Comb:vRegWriteData[15]~1_RESYN1048_BDD1049\,
	datab => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datac => \ALT_INV_Add1~61_sumout\,
	datad => \ALT_INV_Selector17~3_combout\,
	datae => \ALT_INV_R.aluCalc~q\,
	dataf => \ALT_INV_Comb:vRegWriteData[15]~1_RESYN1046_BDD1047\,
	combout => \Comb:vRegWriteData[15]~1_combout\);

-- Location: FF_X80_Y6_N26
\R.regWriteData[15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \R.regWriteData[15]~feeder_combout\,
	asdata => \Comb:vRegWriteData[15]~1_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(15));

-- Location: FF_X73_Y2_N26
\RegFile[31][15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(15),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][15]~q\);

-- Location: LABCELL_X74_Y2_N48
\Mux107~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux107~22_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[24][15]~q\))) # (\R.curInst\(20) & (\RegFile[25][15]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[26][15]~q\))) # (\R.curInst\(20) & (\RegFile[27][15]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[27][15]~q\,
	datab => \ALT_INV_RegFile[25][15]~q\,
	datac => \ALT_INV_RegFile[26][15]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][15]~q\,
	combout => \Mux107~22_combout\);

-- Location: LABCELL_X74_Y2_N24
\Mux107~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux107~9_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux107~22_combout\)))) # (\R.curInst\(22) & ((!\Mux107~22_combout\ & ((\RegFile[28][15]~q\))) # (\Mux107~22_combout\ & (\RegFile[29][15]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux107~22_combout\)))) # (\R.curInst\(22) & ((!\Mux107~22_combout\ & ((\RegFile[30][15]~q\))) # (\Mux107~22_combout\ & (\RegFile[31][15]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][15]~q\,
	datab => \ALT_INV_RegFile[29][15]~q\,
	datac => \ALT_INV_RegFile[30][15]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux107~22_combout\,
	datag => \ALT_INV_RegFile[28][15]~q\,
	combout => \Mux107~9_combout\);

-- Location: LABCELL_X74_Y2_N6
\Mux107~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux107~14_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[8][15]~q\))) # (\R.curInst\(20) & (\RegFile[9][15]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & (\RegFile[10][15]~q\)) # (\R.curInst\(20) & ((\RegFile[11][15]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][15]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[10][15]~q\,
	datad => \ALT_INV_RegFile[11][15]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][15]~q\,
	combout => \Mux107~14_combout\);

-- Location: LABCELL_X74_Y2_N54
\Mux107~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux107~1_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux107~14_combout\)))) # (\R.curInst\(22) & ((!\Mux107~14_combout\ & ((\RegFile[12][15]~q\))) # (\Mux107~14_combout\ & (\RegFile[13][15]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux107~14_combout\)))) # (\R.curInst\(22) & ((!\Mux107~14_combout\ & ((\RegFile[14][15]~q\))) # (\Mux107~14_combout\ & (\RegFile[15][15]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][15]~q\,
	datab => \ALT_INV_RegFile[13][15]~q\,
	datac => \ALT_INV_RegFile[14][15]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux107~14_combout\,
	datag => \ALT_INV_RegFile[12][15]~q\,
	combout => \Mux107~1_combout\);

-- Location: LABCELL_X73_Y1_N51
\Mux107~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux107~18_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & (\RegFile[16][15]~q\)) # (\R.curInst\(20) & ((\RegFile[17][15]~q\)))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & ((\RegFile[18][15]~q\))) # (\R.curInst\(20) & (\RegFile[19][15]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001010101111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[19][15]~q\,
	datac => \ALT_INV_RegFile[18][15]~q\,
	datad => \ALT_INV_RegFile[17][15]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][15]~q\,
	combout => \Mux107~18_combout\);

-- Location: LABCELL_X73_Y1_N12
\Mux107~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux107~5_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux107~18_combout\))))) # (\R.curInst\(22) & (((!\Mux107~18_combout\ & (\RegFile[20][15]~q\)) # (\Mux107~18_combout\ & ((\RegFile[21][15]~q\)))))) ) ) # ( \R.curInst\(21) & ( 
-- (!\R.curInst\(22) & ((((\Mux107~18_combout\))))) # (\R.curInst\(22) & (((!\Mux107~18_combout\ & ((\RegFile[22][15]~q\))) # (\Mux107~18_combout\ & (\RegFile[23][15]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110101010111111111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[23][15]~q\,
	datac => \ALT_INV_RegFile[22][15]~q\,
	datad => \ALT_INV_RegFile[21][15]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux107~18_combout\,
	datag => \ALT_INV_RegFile[20][15]~q\,
	combout => \Mux107~5_combout\);

-- Location: FF_X73_Y3_N37
\RegFile[6][15]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(15),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][15]~DUPLICATE_q\);

-- Location: LABCELL_X71_Y4_N18
\Mux107~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux107~0_combout\ = ( \RegFile[5][15]~q\ & ( \R.curInst\(21) & ( (!\R.curInst\(20) & (\RegFile[6][15]~DUPLICATE_q\)) # (\R.curInst\(20) & ((\RegFile[7][15]~q\))) ) ) ) # ( !\RegFile[5][15]~q\ & ( \R.curInst\(21) & ( (!\R.curInst\(20) & 
-- (\RegFile[6][15]~DUPLICATE_q\)) # (\R.curInst\(20) & ((\RegFile[7][15]~q\))) ) ) ) # ( \RegFile[5][15]~q\ & ( !\R.curInst\(21) & ( (\R.curInst\(20)) # (\RegFile[4][15]~q\) ) ) ) # ( !\RegFile[5][15]~q\ & ( !\R.curInst\(21) & ( (\RegFile[4][15]~q\ & 
-- !\R.curInst\(20)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010100000000010101011111111100110011000011110011001100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[4][15]~q\,
	datab => \ALT_INV_RegFile[6][15]~DUPLICATE_q\,
	datac => \ALT_INV_RegFile[7][15]~q\,
	datad => \ALT_INV_R.curInst\(20),
	datae => \ALT_INV_RegFile[5][15]~q\,
	dataf => \ALT_INV_R.curInst\(21),
	combout => \Mux107~0_combout\);

-- Location: MLABCELL_X72_Y3_N48
\Mux107~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux107~26_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (\RegFile[1][15]~q\ & (\R.curInst\(20)))) # (\R.curInst\(22) & (((\Mux107~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (((\RegFile[2][15]~q\)))) # 
-- (\R.curInst\(20) & (\RegFile[3][15]~q\)))) # (\R.curInst\(22) & ((((\Mux107~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001100000011000100010000110011001111110011111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][15]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[2][15]~q\,
	datad => \ALT_INV_R.curInst\(20),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux107~0_combout\,
	datag => \ALT_INV_RegFile[1][15]~q\,
	combout => \Mux107~26_combout\);

-- Location: LABCELL_X74_Y2_N36
\Mux107~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux107~13_combout\ = ( \Mux107~5_combout\ & ( \Mux107~26_combout\ & ( (!\R.curInst\(23)) # ((!\R.curInst\(24) & ((\Mux107~1_combout\))) # (\R.curInst\(24) & (\Mux107~9_combout\))) ) ) ) # ( !\Mux107~5_combout\ & ( \Mux107~26_combout\ & ( 
-- (!\R.curInst\(23) & (((!\R.curInst\(24))))) # (\R.curInst\(23) & ((!\R.curInst\(24) & ((\Mux107~1_combout\))) # (\R.curInst\(24) & (\Mux107~9_combout\)))) ) ) ) # ( \Mux107~5_combout\ & ( !\Mux107~26_combout\ & ( (!\R.curInst\(23) & (((\R.curInst\(24))))) 
-- # (\R.curInst\(23) & ((!\R.curInst\(24) & ((\Mux107~1_combout\))) # (\R.curInst\(24) & (\Mux107~9_combout\)))) ) ) ) # ( !\Mux107~5_combout\ & ( !\Mux107~26_combout\ & ( (\R.curInst\(23) & ((!\R.curInst\(24) & ((\Mux107~1_combout\))) # (\R.curInst\(24) & 
-- (\Mux107~9_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100010001000000111101110111001111000100011100111111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux107~9_combout\,
	datab => \ALT_INV_R.curInst\(23),
	datac => \ALT_INV_Mux107~1_combout\,
	datad => \ALT_INV_R.curInst\(24),
	datae => \ALT_INV_Mux107~5_combout\,
	dataf => \ALT_INV_Mux107~26_combout\,
	combout => \Mux107~13_combout\);

-- Location: LABCELL_X75_Y6_N27
\NxR.aluData2[15]~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[15]~6_combout\ = ( \Mux107~13_combout\ & ( (!\vAluSrc2~1_combout\) # ((\Mux139~0_combout\ & \Equal4~1_combout\)) ) ) # ( !\Mux107~13_combout\ & ( (\Mux139~0_combout\ & (\vAluSrc2~1_combout\ & \Equal4~1_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000011000000000000001111110000111100111111000011110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Mux139~0_combout\,
	datac => \ALT_INV_vAluSrc2~1_combout\,
	datad => \ALT_INV_Equal4~1_combout\,
	dataf => \ALT_INV_Mux107~13_combout\,
	combout => \NxR.aluData2[15]~6_combout\);

-- Location: FF_X75_Y6_N38
\R.aluData2[15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \NxR.aluData2[15]~6_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData2\(15));

-- Location: LABCELL_X80_Y6_N6
\vAluRes~52\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~52_combout\ = ( !\R.aluCalc~q\ & ( (((\R.aluRes\(15)))) ) ) # ( \R.aluCalc~q\ & ( ((!\Add1~61_sumout\ & (((\R.aluOp.ALUOpSub~q\ & \Add2~61_sumout\)))) # (\Add1~61_sumout\ & (((\R.aluOp.ALUOpSub~q\ & \Add2~61_sumout\)) # (\R.aluOp.ALUOpAdd~q\)))) 
-- # (\Selector17~3_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100001111001101110011011100001111000011110011011111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add1~61_sumout\,
	datab => \ALT_INV_Selector17~3_combout\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datae => \ALT_INV_R.aluCalc~q\,
	dataf => \ALT_INV_Add2~61_sumout\,
	datag => \ALT_INV_R.aluRes\(15),
	combout => \vAluRes~52_combout\);

-- Location: LABCELL_X77_Y5_N30
\Add3~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~1_sumout\ = SUM(( (\R.curInst\(0) & (\R.curInst\(1) & (!\R.curInst\(3) & \Mux154~1_combout\))) ) + ( \R.curPC[0]~DUPLICATE_q\ ) + ( !VCC ))
-- \Add3~2\ = CARRY(( (\R.curInst\(0) & (\R.curInst\(1) & (!\R.curInst\(3) & \Mux154~1_combout\))) ) + ( \R.curPC[0]~DUPLICATE_q\ ) + ( !VCC ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000000000010000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datac => \ALT_INV_R.curInst\(3),
	datad => \ALT_INV_Mux154~1_combout\,
	dataf => \ALT_INV_R.curPC[0]~DUPLICATE_q\,
	cin => GND,
	sumout => \Add3~1_sumout\,
	cout => \Add3~2\);

-- Location: LABCELL_X77_Y5_N33
\Add3~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~5_sumout\ = SUM(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux153~0_combout\)) ) + ( \R.curPC\(1) ) + ( \Add3~2\ ))
-- \Add3~6\ = CARRY(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux153~0_combout\)) ) + ( \R.curPC\(1) ) + ( \Add3~2\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000000100000001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datac => \ALT_INV_Mux153~0_combout\,
	dataf => \ALT_INV_R.curPC\(1),
	cin => \Add3~2\,
	sumout => \Add3~5_sumout\,
	cout => \Add3~6\);

-- Location: LABCELL_X77_Y5_N36
\Add3~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~9_sumout\ = SUM(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux152~0_combout\)) ) + ( \R.curPC\(2) ) + ( \Add3~6\ ))
-- \Add3~10\ = CARRY(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux152~0_combout\)) ) + ( \R.curPC\(2) ) + ( \Add3~6\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000010001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datac => \ALT_INV_R.curPC\(2),
	datad => \ALT_INV_Mux152~0_combout\,
	cin => \Add3~6\,
	sumout => \Add3~9_sumout\,
	cout => \Add3~10\);

-- Location: LABCELL_X77_Y5_N39
\Add3~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~13_sumout\ = SUM(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux151~0_combout\)) ) + ( \R.curPC\(3) ) + ( \Add3~10\ ))
-- \Add3~14\ = CARRY(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux151~0_combout\)) ) + ( \R.curPC\(3) ) + ( \Add3~10\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000000000010001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datad => \ALT_INV_Mux151~0_combout\,
	dataf => \ALT_INV_R.curPC\(3),
	cin => \Add3~10\,
	sumout => \Add3~13_sumout\,
	cout => \Add3~14\);

-- Location: LABCELL_X77_Y5_N42
\Add3~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~17_sumout\ = SUM(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux150~0_combout\)) ) + ( \R.curPC\(4) ) + ( \Add3~14\ ))
-- \Add3~18\ = CARRY(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux150~0_combout\)) ) + ( \R.curPC\(4) ) + ( \Add3~14\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000010001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datac => \ALT_INV_R.curPC\(4),
	datad => \ALT_INV_Mux150~0_combout\,
	cin => \Add3~14\,
	sumout => \Add3~17_sumout\,
	cout => \Add3~18\);

-- Location: LABCELL_X77_Y5_N45
\Add3~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~21_sumout\ = SUM(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux149~1_combout\)) ) + ( \R.curPC\(5) ) + ( \Add3~18\ ))
-- \Add3~22\ = CARRY(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux149~1_combout\)) ) + ( \R.curPC\(5) ) + ( \Add3~18\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000010001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datac => \ALT_INV_R.curPC\(5),
	datad => \ALT_INV_Mux149~1_combout\,
	cin => \Add3~18\,
	sumout => \Add3~21_sumout\,
	cout => \Add3~22\);

-- Location: LABCELL_X77_Y5_N48
\Add3~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~25_sumout\ = SUM(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux148~0_combout\)) ) + ( \R.curPC\(6) ) + ( \Add3~22\ ))
-- \Add3~26\ = CARRY(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux148~0_combout\)) ) + ( \R.curPC\(6) ) + ( \Add3~22\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000000100000001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datac => \ALT_INV_Mux148~0_combout\,
	dataf => \ALT_INV_R.curPC\(6),
	cin => \Add3~22\,
	sumout => \Add3~25_sumout\,
	cout => \Add3~26\);

-- Location: LABCELL_X77_Y5_N51
\Add3~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~29_sumout\ = SUM(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux147~0_combout\)) ) + ( \R.curPC\(7) ) + ( \Add3~26\ ))
-- \Add3~30\ = CARRY(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux147~0_combout\)) ) + ( \R.curPC\(7) ) + ( \Add3~26\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000000100000001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datac => \ALT_INV_Mux147~0_combout\,
	dataf => \ALT_INV_R.curPC\(7),
	cin => \Add3~26\,
	sumout => \Add3~29_sumout\,
	cout => \Add3~30\);

-- Location: LABCELL_X77_Y5_N54
\Add3~33\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~33_sumout\ = SUM(( \R.curPC\(8) ) + ( (\R.curInst\(0) & (\R.curInst\(1) & \Mux146~0_combout\)) ) + ( \Add3~30\ ))
-- \Add3~34\ = CARRY(( \R.curPC\(8) ) + ( (\R.curInst\(0) & (\R.curInst\(1) & \Mux146~0_combout\)) ) + ( \Add3~30\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111101111111000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datac => \ALT_INV_Mux146~0_combout\,
	datad => \ALT_INV_R.curPC\(8),
	cin => \Add3~30\,
	sumout => \Add3~33_sumout\,
	cout => \Add3~34\);

-- Location: LABCELL_X77_Y5_N57
\Add3~37\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~37_sumout\ = SUM(( \R.curPC\(9) ) + ( (\R.curInst\(0) & (\R.curInst\(1) & \Mux145~0_combout\)) ) + ( \Add3~34\ ))
-- \Add3~38\ = CARRY(( \R.curPC\(9) ) + ( (\R.curInst\(0) & (\R.curInst\(1) & \Mux145~0_combout\)) ) + ( \Add3~34\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111101111111000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datac => \ALT_INV_Mux145~0_combout\,
	datad => \ALT_INV_R.curPC\(9),
	cin => \Add3~34\,
	sumout => \Add3~37_sumout\,
	cout => \Add3~38\);

-- Location: LABCELL_X77_Y4_N0
\Add3~41\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~41_sumout\ = SUM(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux144~0_combout\)) ) + ( \R.curPC\(10) ) + ( \Add3~38\ ))
-- \Add3~42\ = CARRY(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux144~0_combout\)) ) + ( \R.curPC\(10) ) + ( \Add3~38\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000000000010001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datad => \ALT_INV_Mux144~0_combout\,
	dataf => \ALT_INV_R.curPC\(10),
	cin => \Add3~38\,
	sumout => \Add3~41_sumout\,
	cout => \Add3~42\);

-- Location: LABCELL_X77_Y4_N3
\Add3~45\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~45_sumout\ = SUM(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux143~1_combout\)) ) + ( \R.curPC\(11) ) + ( \Add3~42\ ))
-- \Add3~46\ = CARRY(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux143~1_combout\)) ) + ( \R.curPC\(11) ) + ( \Add3~42\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000000100000001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datac => \ALT_INV_Mux143~1_combout\,
	dataf => \ALT_INV_R.curPC\(11),
	cin => \Add3~42\,
	sumout => \Add3~45_sumout\,
	cout => \Add3~46\);

-- Location: LABCELL_X77_Y4_N6
\Add3~49\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~49_sumout\ = SUM(( \R.curPC\(12) ) + ( (\R.curInst\(0) & (\R.curInst\(1) & \Mux142~0_combout\)) ) + ( \Add3~46\ ))
-- \Add3~50\ = CARRY(( \R.curPC\(12) ) + ( (\R.curInst\(0) & (\R.curInst\(1) & \Mux142~0_combout\)) ) + ( \Add3~46\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111101111111000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datac => \ALT_INV_Mux142~0_combout\,
	datad => \ALT_INV_R.curPC\(12),
	cin => \Add3~46\,
	sumout => \Add3~49_sumout\,
	cout => \Add3~50\);

-- Location: LABCELL_X77_Y4_N9
\Add3~53\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~53_sumout\ = SUM(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux141~0_combout\)) ) + ( \R.curPC\(13) ) + ( \Add3~50\ ))
-- \Add3~54\ = CARRY(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux141~0_combout\)) ) + ( \R.curPC\(13) ) + ( \Add3~50\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000010001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datac => \ALT_INV_R.curPC\(13),
	datad => \ALT_INV_Mux141~0_combout\,
	cin => \Add3~50\,
	sumout => \Add3~53_sumout\,
	cout => \Add3~54\);

-- Location: LABCELL_X77_Y4_N12
\Add3~57\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~57_sumout\ = SUM(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux140~0_combout\)) ) + ( \R.curPC\(14) ) + ( \Add3~54\ ))
-- \Add3~58\ = CARRY(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux140~0_combout\)) ) + ( \R.curPC\(14) ) + ( \Add3~54\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000000100000001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datac => \ALT_INV_Mux140~0_combout\,
	dataf => \ALT_INV_R.curPC\(14),
	cin => \Add3~54\,
	sumout => \Add3~57_sumout\,
	cout => \Add3~58\);

-- Location: LABCELL_X77_Y4_N15
\Add3~61\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~61_sumout\ = SUM(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux139~0_combout\)) ) + ( \R.curPC\(15) ) + ( \Add3~58\ ))
-- \Add3~62\ = CARRY(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux139~0_combout\)) ) + ( \R.curPC\(15) ) + ( \Add3~58\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000000000000101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datac => \ALT_INV_R.curInst\(1),
	datad => \ALT_INV_Mux139~0_combout\,
	dataf => \ALT_INV_R.curPC\(15),
	cin => \Add3~58\,
	sumout => \Add3~61_sumout\,
	cout => \Add3~62\);

-- Location: LABCELL_X80_Y6_N54
\Comb:vJumpAdr[15]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[15]~0_combout\ = ( \Add3~61_sumout\ & ( (!\Equal4~2_combout\) # (\vAluRes~52_combout\) ) ) # ( !\Add3~61_sumout\ & ( (\vAluRes~52_combout\ & \Equal4~2_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110011000000000011001111111111001100111111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_vAluRes~52_combout\,
	datad => \ALT_INV_Equal4~2_combout\,
	dataf => \ALT_INV_Add3~61_sumout\,
	combout => \Comb:vJumpAdr[15]~0_combout\);

-- Location: MLABCELL_X78_Y1_N24
\Mux44~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux44~0_combout\ = ( \R.curInst\(5) & ( (\R.curInst\(4) & (\R.curInst\(0) & \R.curInst\(6))) ) ) # ( !\R.curInst\(5) & ( (!\R.curInst\(4) & (\R.curInst\(0) & !\R.curInst\(6))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000110000000000000011000000000000000000000000110000000000000011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.curInst\(4),
	datac => \ALT_INV_R.curInst\(0),
	datad => \ALT_INV_R.curInst\(6),
	dataf => \ALT_INV_R.curInst\(5),
	combout => \Mux44~0_combout\);

-- Location: MLABCELL_X78_Y1_N39
\NxR~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR~10_combout\ = ( \R.ctrlState.Calc~q\ & ( \Mux44~0_combout\ & ( (\R.curInst\(1) & \Mux53~0_combout\) ) ) ) # ( !\R.ctrlState.Calc~q\ & ( \Mux44~0_combout\ & ( \R.ctrlState.CheckJump~q\ ) ) ) # ( !\R.ctrlState.Calc~q\ & ( !\Mux44~0_combout\ & ( 
-- \R.ctrlState.CheckJump~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110011000000000000000000110011001100110000010100000101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(1),
	datab => \ALT_INV_R.ctrlState.CheckJump~q\,
	datac => \ALT_INV_Mux53~0_combout\,
	datae => \ALT_INV_R.ctrlState.Calc~q\,
	dataf => \ALT_INV_Mux44~0_combout\,
	combout => \NxR~10_combout\);

-- Location: MLABCELL_X78_Y1_N21
\NxR~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR~9_combout\ = ( \R.curInst\(5) & ( (\R.curInst\(6) & ((!\R.curInst\(4)) # (!\Mux0~0_combout\))) ) ) # ( !\R.curInst\(5) & ( (!\R.curInst\(6) & !\R.curInst\(4)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000100010001000100010001000100001010101010001000101010101000100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(6),
	datab => \ALT_INV_R.curInst\(4),
	datad => \ALT_INV_Mux0~0_combout\,
	dataf => \ALT_INV_R.curInst\(5),
	combout => \NxR~9_combout\);

-- Location: MLABCELL_X78_Y1_N12
\NxR~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR~11_combout\ = ( \Mux53~1_combout\ & ( (!\R.ctrlState.ReadReg~q\ & (\NxR~10_combout\)) # (\R.ctrlState.ReadReg~q\ & ((!\NxR~9_combout\))) ) ) # ( !\Mux53~1_combout\ & ( (\NxR~10_combout\) # (\R.ctrlState.ReadReg~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0111011101110111011101110111011101110010011100100111001001110010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.ctrlState.ReadReg~q\,
	datab => \ALT_INV_NxR~10_combout\,
	datac => \ALT_INV_NxR~9_combout\,
	dataf => \ALT_INV_Mux53~1_combout\,
	combout => \NxR~11_combout\);

-- Location: FF_X78_Y1_N13
\R.incPC\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR~11_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sclr => \R.ctrlState.Fetch~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.incPC~q\);

-- Location: MLABCELL_X78_Y4_N33
\NxR.curPC[31]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.curPC[31]~0_combout\ = (\R.incPC~q\) # (\R.jumpToAdr~q\)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111111111111000011111111111100001111111111110000111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.jumpToAdr~q\,
	datad => \ALT_INV_R.incPC~q\,
	combout => \NxR.curPC[31]~0_combout\);

-- Location: FF_X80_Y6_N55
\R.curPC[15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[15]~0_combout\,
	asdata => \Add0~53_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(15));

-- Location: LABCELL_X81_Y6_N45
\Add0~61\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~61_sumout\ = SUM(( \R.curPC\(17) ) + ( GND ) + ( \Add0~58\ ))
-- \Add0~62\ = CARRY(( \R.curPC\(17) ) + ( GND ) + ( \Add0~58\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.curPC\(17),
	cin => \Add0~58\,
	sumout => \Add0~61_sumout\,
	cout => \Add0~62\);

-- Location: MLABCELL_X78_Y3_N3
\R.regWriteData[17]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.regWriteData[17]~feeder_combout\ = ( \Add0~61_sumout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_Add0~61_sumout\,
	combout => \R.regWriteData[17]~feeder_combout\);

-- Location: MLABCELL_X78_Y3_N33
\Comb:vRegWriteData[17]~1_RESYN1124\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[17]~1_RESYN1124_BDD1125\ = (\R.aluCalc~q\ & !\R.memToReg~q\)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101000001010000010100000101000001010000010100000101000001010000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_R.memToReg~q\,
	combout => \Comb:vRegWriteData[17]~1_RESYN1124_BDD1125\);

-- Location: IOIBUF_X58_Y0_N92
\avm_d_readdata[9]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(9),
	o => \avm_d_readdata[9]~input_o\);

-- Location: LABCELL_X79_Y2_N30
\Comb:vRegWriteData[17]~1_RESYN1120\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[17]~1_RESYN1120_BDD1121\ = ( \avm_d_readdata[23]~input_o\ & ( \avm_d_readdata[9]~input_o\ & ( (!\R.curInst\(14) & ((!\R.curInst\(12) & ((\R.curInst\(13)) # (\avm_d_readdata[31]~input_o\))) # (\R.curInst\(12) & ((!\R.curInst\(13)))))) ) 
-- ) ) # ( !\avm_d_readdata[23]~input_o\ & ( \avm_d_readdata[9]~input_o\ & ( (!\R.curInst\(12) & (!\R.curInst\(14) & ((\R.curInst\(13)) # (\avm_d_readdata[31]~input_o\)))) ) ) ) # ( \avm_d_readdata[23]~input_o\ & ( !\avm_d_readdata[9]~input_o\ & ( 
-- (!\R.curInst\(13) & (!\R.curInst\(14) & ((\avm_d_readdata[31]~input_o\) # (\R.curInst\(12))))) ) ) ) # ( !\avm_d_readdata[23]~input_o\ & ( !\avm_d_readdata[9]~input_o\ & ( (!\R.curInst\(12) & (\avm_d_readdata[31]~input_o\ & (!\R.curInst\(13) & 
-- !\R.curInst\(14)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010000000000000011100000000000000101010000000000111101000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(12),
	datab => \ALT_INV_avm_d_readdata[31]~input_o\,
	datac => \ALT_INV_R.curInst\(13),
	datad => \ALT_INV_R.curInst\(14),
	datae => \ALT_INV_avm_d_readdata[23]~input_o\,
	dataf => \ALT_INV_avm_d_readdata[9]~input_o\,
	combout => \Comb:vRegWriteData[17]~1_RESYN1120_BDD1121\);

-- Location: MLABCELL_X78_Y3_N6
\Comb:vRegWriteData[17]~1_RESYN1122\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[17]~1_RESYN1122_BDD1123\ = ( \R.aluOp.ALUOpSub~q\ & ( \Comb:vRegWriteData[17]~1_RESYN1120_BDD1121\ & ( ((!\R.aluCalc~q\ & (\R.aluRes\(17))) # (\R.aluCalc~q\ & ((\Add2~69_sumout\)))) # (\R.memToReg~q\) ) ) ) # ( !\R.aluOp.ALUOpSub~q\ & 
-- ( \Comb:vRegWriteData[17]~1_RESYN1120_BDD1121\ & ( ((\R.aluRes\(17) & !\R.aluCalc~q\)) # (\R.memToReg~q\) ) ) ) # ( \R.aluOp.ALUOpSub~q\ & ( !\Comb:vRegWriteData[17]~1_RESYN1120_BDD1121\ & ( (!\R.memToReg~q\ & ((!\R.aluCalc~q\ & (\R.aluRes\(17))) # 
-- (\R.aluCalc~q\ & ((\Add2~69_sumout\))))) ) ) ) # ( !\R.aluOp.ALUOpSub~q\ & ( !\Comb:vRegWriteData[17]~1_RESYN1120_BDD1121\ & ( (\R.aluRes\(17) & (!\R.aluCalc~q\ & !\R.memToReg~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100010000000000010001110000000001000100111111110100011111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluRes\(17),
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_Add2~69_sumout\,
	datad => \ALT_INV_R.memToReg~q\,
	datae => \ALT_INV_R.aluOp.ALUOpSub~q\,
	dataf => \ALT_INV_Comb:vRegWriteData[17]~1_RESYN1120_BDD1121\,
	combout => \Comb:vRegWriteData[17]~1_RESYN1122_BDD1123\);

-- Location: MLABCELL_X78_Y3_N18
\Comb:vRegWriteData[17]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[17]~1_combout\ = ( \Selector15~0_combout\ & ( \Comb:vRegWriteData[17]~1_RESYN1122_BDD1123\ ) ) # ( !\Selector15~0_combout\ & ( \Comb:vRegWriteData[17]~1_RESYN1122_BDD1123\ ) ) # ( \Selector15~0_combout\ & ( 
-- !\Comb:vRegWriteData[17]~1_RESYN1122_BDD1123\ & ( \Comb:vRegWriteData[17]~1_RESYN1124_BDD1125\ ) ) ) # ( !\Selector15~0_combout\ & ( !\Comb:vRegWriteData[17]~1_RESYN1122_BDD1123\ & ( (\Comb:vRegWriteData[17]~1_RESYN1124_BDD1125\ & 
-- ((!\Selector15~4_combout\) # ((\R.aluOp.ALUOpAdd~q\ & \Add1~69_sumout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000110000001101000011110000111111111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datab => \ALT_INV_Selector15~4_combout\,
	datac => \ALT_INV_Comb:vRegWriteData[17]~1_RESYN1124_BDD1125\,
	datad => \ALT_INV_Add1~69_sumout\,
	datae => \ALT_INV_Selector15~0_combout\,
	dataf => \ALT_INV_Comb:vRegWriteData[17]~1_RESYN1122_BDD1123\,
	combout => \Comb:vRegWriteData[17]~1_combout\);

-- Location: FF_X78_Y3_N5
\R.regWriteData[17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \R.regWriteData[17]~feeder_combout\,
	asdata => \Comb:vRegWriteData[17]~1_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(17));

-- Location: FF_X62_Y5_N38
\RegFile[13][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(17),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][17]~q\);

-- Location: LABCELL_X64_Y3_N6
\Mux105~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux105~14_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[8][17]~q\))) # (\R.curInst\(20) & (\RegFile[9][17]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[10][17]~q\))) # (\R.curInst\(20) & (\RegFile[11][17]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[11][17]~q\,
	datab => \ALT_INV_RegFile[9][17]~q\,
	datac => \ALT_INV_RegFile[10][17]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][17]~q\,
	combout => \Mux105~14_combout\);

-- Location: LABCELL_X62_Y5_N36
\Mux105~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux105~1_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux105~14_combout\))))) # (\R.curInst\(22) & (((!\Mux105~14_combout\ & ((\RegFile[12][17]~q\))) # (\Mux105~14_combout\ & (\RegFile[13][17]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux105~14_combout\)))) # (\R.curInst\(22) & ((!\Mux105~14_combout\ & (\RegFile[14][17]~q\)) # (\Mux105~14_combout\ & ((\RegFile[15][17]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][17]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[14][17]~q\,
	datad => \ALT_INV_RegFile[15][17]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux105~14_combout\,
	datag => \ALT_INV_RegFile[12][17]~q\,
	combout => \Mux105~1_combout\);

-- Location: LABCELL_X63_Y5_N54
\Mux105~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux105~18_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[16][17]~q\))) # (\R.curInst\(20) & (\RegFile[17][17]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & (\RegFile[18][17]~q\)) # (\R.curInst\(20) & ((\RegFile[19][17]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[17][17]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[18][17]~q\,
	datad => \ALT_INV_RegFile[19][17]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][17]~q\,
	combout => \Mux105~18_combout\);

-- Location: LABCELL_X63_Y5_N48
\Mux105~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux105~5_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux105~18_combout\)))) # (\R.curInst\(22) & ((!\Mux105~18_combout\ & ((\RegFile[20][17]~q\))) # (\Mux105~18_combout\ & (\RegFile[21][17]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux105~18_combout\)))) # (\R.curInst\(22) & ((!\Mux105~18_combout\ & ((\RegFile[22][17]~q\))) # (\Mux105~18_combout\ & (\RegFile[23][17]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][17]~q\,
	datab => \ALT_INV_RegFile[23][17]~q\,
	datac => \ALT_INV_RegFile[22][17]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux105~18_combout\,
	datag => \ALT_INV_RegFile[20][17]~q\,
	combout => \Mux105~5_combout\);

-- Location: LABCELL_X61_Y2_N30
\Mux105~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux105~0_combout\ = ( \RegFile[5][17]~q\ & ( \R.curInst\(20) & ( (!\R.curInst\(21)) # (\RegFile[7][17]~q\) ) ) ) # ( !\RegFile[5][17]~q\ & ( \R.curInst\(20) & ( (\RegFile[7][17]~q\ & \R.curInst\(21)) ) ) ) # ( \RegFile[5][17]~q\ & ( !\R.curInst\(20) & ( 
-- (!\R.curInst\(21) & ((\RegFile[4][17]~q\))) # (\R.curInst\(21) & (\RegFile[6][17]~q\)) ) ) ) # ( !\RegFile[5][17]~q\ & ( !\R.curInst\(20) & ( (!\R.curInst\(21) & ((\RegFile[4][17]~q\))) # (\R.curInst\(21) & (\RegFile[6][17]~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001101010101001100110101010100000000000011111111111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[6][17]~q\,
	datab => \ALT_INV_RegFile[4][17]~q\,
	datac => \ALT_INV_RegFile[7][17]~q\,
	datad => \ALT_INV_R.curInst\(21),
	datae => \ALT_INV_RegFile[5][17]~q\,
	dataf => \ALT_INV_R.curInst\(20),
	combout => \Mux105~0_combout\);

-- Location: FF_X61_Y5_N23
\RegFile[1][17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(17),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][17]~q\);

-- Location: LABCELL_X61_Y5_N6
\Mux105~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux105~26_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((\RegFile[1][17]~q\ & (\R.curInst\(20)))))) # (\R.curInst\(22) & ((((\Mux105~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (((\RegFile[2][17]~q\)))) 
-- # (\R.curInst\(20) & (\RegFile[3][17]~q\)))) # (\R.curInst\(22) & ((((\Mux105~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001010000010100010001001010101010111110101111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[3][17]~q\,
	datac => \ALT_INV_RegFile[2][17]~q\,
	datad => \ALT_INV_R.curInst\(20),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux105~0_combout\,
	datag => \ALT_INV_RegFile[1][17]~q\,
	combout => \Mux105~26_combout\);

-- Location: LABCELL_X62_Y4_N36
\Mux105~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux105~22_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[24][17]~q\))) # (\R.curInst\(20) & (\RegFile[25][17]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[26][17]~q\))) # (\R.curInst\(20) & (\RegFile[27][17]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[25][17]~q\,
	datab => \ALT_INV_RegFile[27][17]~q\,
	datac => \ALT_INV_RegFile[26][17]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][17]~q\,
	combout => \Mux105~22_combout\);

-- Location: LABCELL_X62_Y5_N42
\Mux105~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux105~9_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux105~22_combout\)))) # (\R.curInst\(22) & ((!\Mux105~22_combout\ & ((\RegFile[28][17]~q\))) # (\Mux105~22_combout\ & (\RegFile[29][17]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux105~22_combout\)))) # (\R.curInst\(22) & ((!\Mux105~22_combout\ & ((\RegFile[30][17]~q\))) # (\Mux105~22_combout\ & (\RegFile[31][17]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[29][17]~q\,
	datab => \ALT_INV_RegFile[31][17]~q\,
	datac => \ALT_INV_RegFile[30][17]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux105~22_combout\,
	datag => \ALT_INV_RegFile[28][17]~q\,
	combout => \Mux105~9_combout\);

-- Location: LABCELL_X62_Y5_N48
\Mux105~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux105~13_combout\ = ( \Mux105~26_combout\ & ( \Mux105~9_combout\ & ( (!\R.curInst\(24) & (((!\R.curInst\(23))) # (\Mux105~1_combout\))) # (\R.curInst\(24) & (((\R.curInst\(23)) # (\Mux105~5_combout\)))) ) ) ) # ( !\Mux105~26_combout\ & ( 
-- \Mux105~9_combout\ & ( (!\R.curInst\(24) & (\Mux105~1_combout\ & ((\R.curInst\(23))))) # (\R.curInst\(24) & (((\R.curInst\(23)) # (\Mux105~5_combout\)))) ) ) ) # ( \Mux105~26_combout\ & ( !\Mux105~9_combout\ & ( (!\R.curInst\(24) & (((!\R.curInst\(23))) # 
-- (\Mux105~1_combout\))) # (\R.curInst\(24) & (((\Mux105~5_combout\ & !\R.curInst\(23))))) ) ) ) # ( !\Mux105~26_combout\ & ( !\Mux105~9_combout\ & ( (!\R.curInst\(24) & (\Mux105~1_combout\ & ((\R.curInst\(23))))) # (\R.curInst\(24) & (((\Mux105~5_combout\ 
-- & !\R.curInst\(23))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001101010000111100110101000000000011010111111111001101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux105~1_combout\,
	datab => \ALT_INV_Mux105~5_combout\,
	datac => \ALT_INV_R.curInst\(24),
	datad => \ALT_INV_R.curInst\(23),
	datae => \ALT_INV_Mux105~26_combout\,
	dataf => \ALT_INV_Mux105~9_combout\,
	combout => \Mux105~13_combout\);

-- Location: MLABCELL_X72_Y5_N3
\NxR.aluData2[17]~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[17]~4_combout\ = ( \Mux105~13_combout\ & ( (!\vAluSrc2~1_combout\) # ((\Mux137~0_combout\ & \Equal4~1_combout\)) ) ) # ( !\Mux105~13_combout\ & ( (\Mux137~0_combout\ & (\Equal4~1_combout\ & \vAluSrc2~1_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000011000000000000001111111111000000111111111100000011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Mux137~0_combout\,
	datac => \ALT_INV_Equal4~1_combout\,
	datad => \ALT_INV_vAluSrc2~1_combout\,
	dataf => \ALT_INV_Mux105~13_combout\,
	combout => \NxR.aluData2[17]~4_combout\);

-- Location: FF_X72_Y5_N34
\Add2~65_OTERM703_NEW_REG806\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \NxR.aluData2[17]~4_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Add2~65_OTERM703_OTERM807\);

-- Location: MLABCELL_X78_Y3_N54
\Selector15~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector15~5_combout\ = ( \Add1~69_sumout\ & ( \Selector15~4_combout\ & ( (((\Add2~69_sumout\ & \R.aluOp.ALUOpSub~q\)) # (\Selector15~0_combout\)) # (\R.aluOp.ALUOpAdd~q\) ) ) ) # ( !\Add1~69_sumout\ & ( \Selector15~4_combout\ & ( ((\Add2~69_sumout\ & 
-- \R.aluOp.ALUOpSub~q\)) # (\Selector15~0_combout\) ) ) ) # ( \Add1~69_sumout\ & ( !\Selector15~4_combout\ ) ) # ( !\Add1~69_sumout\ & ( !\Selector15~4_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111111111111111111100010001111111110001111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add2~69_sumout\,
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_Selector15~0_combout\,
	datae => \ALT_INV_Add1~69_sumout\,
	dataf => \ALT_INV_Selector15~4_combout\,
	combout => \Selector15~5_combout\);

-- Location: LABCELL_X77_Y4_N18
\Add3~65\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~65_sumout\ = SUM(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux138~0_combout\)) ) + ( \R.curPC\(16) ) + ( \Add3~62\ ))
-- \Add3~66\ = CARRY(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux138~0_combout\)) ) + ( \R.curPC\(16) ) + ( \Add3~62\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000000000010001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datad => \ALT_INV_Mux138~0_combout\,
	dataf => \ALT_INV_R.curPC\(16),
	cin => \Add3~62\,
	sumout => \Add3~65_sumout\,
	cout => \Add3~66\);

-- Location: LABCELL_X77_Y4_N21
\Add3~69\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~69_sumout\ = SUM(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux137~0_combout\)) ) + ( \R.curPC\(17) ) + ( \Add3~66\ ))
-- \Add3~70\ = CARRY(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux137~0_combout\)) ) + ( \R.curPC\(17) ) + ( \Add3~66\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000000000000101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datac => \ALT_INV_R.curInst\(1),
	datad => \ALT_INV_Mux137~0_combout\,
	dataf => \ALT_INV_R.curPC\(17),
	cin => \Add3~66\,
	sumout => \Add3~69_sumout\,
	cout => \Add3~70\);

-- Location: MLABCELL_X78_Y3_N30
\Comb:vJumpAdr[17]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[17]~0_combout\ = ( \Add3~69_sumout\ & ( (!\Equal4~2_combout\) # ((!\R.aluCalc~q\ & ((\R.aluRes\(17)))) # (\R.aluCalc~q\ & (\Selector15~5_combout\))) ) ) # ( !\Add3~69_sumout\ & ( (\Equal4~2_combout\ & ((!\R.aluCalc~q\ & ((\R.aluRes\(17)))) 
-- # (\R.aluCalc~q\ & (\Selector15~5_combout\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000100100011000000010010001111001101111011111100110111101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluCalc~q\,
	datab => \ALT_INV_Equal4~2_combout\,
	datac => \ALT_INV_Selector15~5_combout\,
	datad => \ALT_INV_R.aluRes\(17),
	dataf => \ALT_INV_Add3~69_sumout\,
	combout => \Comb:vJumpAdr[17]~0_combout\);

-- Location: FF_X78_Y3_N31
\R.curPC[17]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[17]~0_combout\,
	asdata => \Add0~61_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(17));

-- Location: LABCELL_X81_Y6_N48
\Add0~65\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~65_sumout\ = SUM(( \R.curPC\(18) ) + ( GND ) + ( \Add0~62\ ))
-- \Add0~66\ = CARRY(( \R.curPC\(18) ) + ( GND ) + ( \Add0~62\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.curPC\(18),
	cin => \Add0~62\,
	sumout => \Add0~65_sumout\,
	cout => \Add0~66\);

-- Location: LABCELL_X79_Y3_N45
\R.regWriteData[18]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.regWriteData[18]~feeder_combout\ = ( \Add0~65_sumout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_Add0~65_sumout\,
	combout => \R.regWriteData[18]~feeder_combout\);

-- Location: IOIBUF_X34_Y0_N92
\avm_d_readdata[10]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(10),
	o => \avm_d_readdata[10]~input_o\);

-- Location: LABCELL_X79_Y2_N21
\Comb:vRegWriteData[18]~1_RESYN1736\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[18]~1_RESYN1736_BDD1737\ = ( \R.curInst\(12) & ( (\avm_d_readdata[23]~input_o\ & !\R.curInst\(13)) ) ) # ( !\R.curInst\(12) & ( (!\R.curInst\(13) & (\avm_d_readdata[31]~input_o\)) # (\R.curInst\(13) & ((\avm_d_readdata[10]~input_o\))) 
-- ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100001111001100110000111101010101000000000101010100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_avm_d_readdata[23]~input_o\,
	datab => \ALT_INV_avm_d_readdata[31]~input_o\,
	datac => \ALT_INV_avm_d_readdata[10]~input_o\,
	datad => \ALT_INV_R.curInst\(13),
	dataf => \ALT_INV_R.curInst\(12),
	combout => \Comb:vRegWriteData[18]~1_RESYN1736_BDD1737\);

-- Location: LABCELL_X80_Y3_N18
\Comb:vRegWriteData[18]~1_RESYN1738\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[18]~1_RESYN1738_BDD1739\ = ( \Comb:vRegWriteData[24]~1_combout\ & ( \Comb:vRegWriteData[18]~1_RESYN1736_BDD1737\ ) ) # ( !\Comb:vRegWriteData[24]~1_combout\ & ( \Comb:vRegWriteData[18]~1_RESYN1736_BDD1737\ & ( (!\R.aluCalc~q\ & 
-- (\R.aluRes\(18) & !\R.memToReg~q\)) ) ) ) # ( \Comb:vRegWriteData[24]~1_combout\ & ( !\Comb:vRegWriteData[18]~1_RESYN1736_BDD1737\ & ( (!\R.aluCalc~q\ & (\R.aluRes\(18) & !\R.memToReg~q\)) ) ) ) # ( !\Comb:vRegWriteData[24]~1_combout\ & ( 
-- !\Comb:vRegWriteData[18]~1_RESYN1736_BDD1737\ & ( (!\R.aluCalc~q\ & (\R.aluRes\(18) & !\R.memToReg~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010000000100000001000000010000000100000001000001111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluCalc~q\,
	datab => \ALT_INV_R.aluRes\(18),
	datac => \ALT_INV_R.memToReg~q\,
	datae => \ALT_INV_Comb:vRegWriteData[24]~1_combout\,
	dataf => \ALT_INV_Comb:vRegWriteData[18]~1_RESYN1736_BDD1737\,
	combout => \Comb:vRegWriteData[18]~1_RESYN1738_BDD1739\);

-- Location: LABCELL_X79_Y3_N30
\Comb:vRegWriteData[18]~1_RESYN1740\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[18]~1_RESYN1740_BDD1741\ = ( \R.memToReg~q\ & ( \Comb:vRegWriteData[18]~1_RESYN1738_BDD1739\ ) ) # ( !\R.memToReg~q\ & ( \Comb:vRegWriteData[18]~1_RESYN1738_BDD1739\ ) ) # ( !\R.memToReg~q\ & ( 
-- !\Comb:vRegWriteData[18]~1_RESYN1738_BDD1739\ & ( (\R.aluCalc~q\ & ((!\Selector14~2_combout\) # ((\Add2~73_sumout\ & \R.aluOp.ALUOpSub~q\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010100000001000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluCalc~q\,
	datab => \ALT_INV_Add2~73_sumout\,
	datac => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datad => \ALT_INV_Selector14~2_combout\,
	datae => \ALT_INV_R.memToReg~q\,
	dataf => \ALT_INV_Comb:vRegWriteData[18]~1_RESYN1738_BDD1739\,
	combout => \Comb:vRegWriteData[18]~1_RESYN1740_BDD1741\);

-- Location: LABCELL_X79_Y3_N36
\Comb:vRegWriteData[18]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[18]~1_combout\ = ( \Add1~73_sumout\ & ( \Comb:vRegWriteData[18]~1_RESYN1740_BDD1741\ ) ) # ( !\Add1~73_sumout\ & ( \Comb:vRegWriteData[18]~1_RESYN1740_BDD1741\ ) ) # ( \Add1~73_sumout\ & ( !\Comb:vRegWriteData[18]~1_RESYN1740_BDD1741\ 
-- & ( (\R.aluCalc~q\ & (!\R.memToReg~q\ & ((\Selector14~4_combout\) # (\R.aluOp.ALUOpAdd~q\)))) ) ) ) # ( !\Add1~73_sumout\ & ( !\Comb:vRegWriteData[18]~1_RESYN1740_BDD1741\ & ( (\R.aluCalc~q\ & (!\R.memToReg~q\ & \Selector14~4_combout\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001000100000001000100010011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluCalc~q\,
	datab => \ALT_INV_R.memToReg~q\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_Selector14~4_combout\,
	datae => \ALT_INV_Add1~73_sumout\,
	dataf => \ALT_INV_Comb:vRegWriteData[18]~1_RESYN1740_BDD1741\,
	combout => \Comb:vRegWriteData[18]~1_combout\);

-- Location: FF_X79_Y3_N47
\R.regWriteData[18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \R.regWriteData[18]~feeder_combout\,
	asdata => \Comb:vRegWriteData[18]~1_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(18));

-- Location: FF_X68_Y7_N32
\RegFile[21][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(18),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][18]~q\);

-- Location: LABCELL_X64_Y4_N24
\Mux72~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux72~18_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & (\RegFile[16][18]~q\)) # (\R.curInst\(15) & ((\RegFile[17][18]~q\)))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & ((\RegFile[18][18]~q\))) # (\R.curInst\(15) & (\RegFile[19][18]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001010101111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[19][18]~q\,
	datac => \ALT_INV_RegFile[18][18]~q\,
	datad => \ALT_INV_RegFile[17][18]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][18]~q\,
	combout => \Mux72~18_combout\);

-- Location: LABCELL_X64_Y4_N12
\Mux72~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux72~5_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux72~18_combout\))))) # (\R.curInst\(17) & (((!\Mux72~18_combout\ & ((\RegFile[20][18]~q\))) # (\Mux72~18_combout\ & (\RegFile[21][18]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux72~18_combout\)))) # (\R.curInst\(17) & ((!\Mux72~18_combout\ & (\RegFile[22][18]~q\)) # (\Mux72~18_combout\ & ((\RegFile[23][18]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][18]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[22][18]~q\,
	datad => \ALT_INV_RegFile[23][18]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux72~18_combout\,
	datag => \ALT_INV_RegFile[20][18]~q\,
	combout => \Mux72~5_combout\);

-- Location: FF_X67_Y5_N37
\RegFile[4][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(18),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][18]~q\);

-- Location: FF_X68_Y4_N38
\RegFile[6][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[6][18]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][18]~q\);

-- Location: LABCELL_X68_Y4_N18
\Mux72~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux72~0_combout\ = ( \RegFile[7][18]~q\ & ( \R.curInst\(15) & ( (\RegFile[5][18]~q\) # (\R.curInst\(16)) ) ) ) # ( !\RegFile[7][18]~q\ & ( \R.curInst\(15) & ( (!\R.curInst\(16) & \RegFile[5][18]~q\) ) ) ) # ( \RegFile[7][18]~q\ & ( !\R.curInst\(15) & ( 
-- (!\R.curInst\(16) & (\RegFile[4][18]~q\)) # (\R.curInst\(16) & ((\RegFile[6][18]~q\))) ) ) ) # ( !\RegFile[7][18]~q\ & ( !\R.curInst\(15) & ( (!\R.curInst\(16) & (\RegFile[4][18]~q\)) # (\R.curInst\(16) & ((\RegFile[6][18]~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100011101000111010001110100011100000000110011000011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[4][18]~q\,
	datab => \ALT_INV_R.curInst\(16),
	datac => \ALT_INV_RegFile[6][18]~q\,
	datad => \ALT_INV_RegFile[5][18]~q\,
	datae => \ALT_INV_RegFile[7][18]~q\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux72~0_combout\);

-- Location: LABCELL_X68_Y4_N6
\Mux72~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux72~26_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((\RegFile[1][18]~q\ & (\R.curInst\(15)))))) # (\R.curInst\(17) & ((((\Mux72~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & ((!\R.curInst\(15) & (((\RegFile[2][18]~q\)))) # 
-- (\R.curInst\(15) & (\RegFile[3][18]~q\)))) # (\R.curInst\(17) & ((((\Mux72~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001010000010100010001001010101010111110101111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[3][18]~q\,
	datac => \ALT_INV_RegFile[2][18]~q\,
	datad => \ALT_INV_R.curInst\(15),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux72~0_combout\,
	datag => \ALT_INV_RegFile[1][18]~q\,
	combout => \Mux72~26_combout\);

-- Location: FF_X62_Y6_N32
\RegFile[30][18]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[30][18]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][18]~DUPLICATE_q\);

-- Location: LABCELL_X62_Y4_N48
\Mux72~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux72~22_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & (\RegFile[24][18]~q\)) # (\R.curInst\(15) & ((\RegFile[25][18]~q\)))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & ((\RegFile[26][18]~q\))) # (\R.curInst\(15) & (\RegFile[27][18]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001010101111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[27][18]~q\,
	datac => \ALT_INV_RegFile[26][18]~q\,
	datad => \ALT_INV_RegFile[25][18]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][18]~q\,
	combout => \Mux72~22_combout\);

-- Location: LABCELL_X62_Y4_N12
\Mux72~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux72~9_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux72~22_combout\))))) # (\R.curInst\(17) & (((!\Mux72~22_combout\ & ((\RegFile[28][18]~q\))) # (\Mux72~22_combout\ & (\RegFile[29][18]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- (!\R.curInst\(17) & ((((\Mux72~22_combout\))))) # (\R.curInst\(17) & (((!\Mux72~22_combout\ & (\RegFile[30][18]~DUPLICATE_q\)) # (\Mux72~22_combout\ & ((\RegFile[31][18]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110111011101110111010101011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[29][18]~q\,
	datac => \ALT_INV_RegFile[30][18]~DUPLICATE_q\,
	datad => \ALT_INV_RegFile[31][18]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux72~22_combout\,
	datag => \ALT_INV_RegFile[28][18]~q\,
	combout => \Mux72~9_combout\);

-- Location: FF_X65_Y3_N56
\RegFile[10][18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[10][18]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][18]~q\);

-- Location: MLABCELL_X65_Y3_N24
\Mux72~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux72~14_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[8][18]~q\))) # (\R.curInst\(15) & (\RegFile[9][18]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & (\RegFile[10][18]~q\)) # (\R.curInst\(15) & ((\RegFile[11][18]~q\))))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][18]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[10][18]~q\,
	datad => \ALT_INV_RegFile[11][18]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][18]~q\,
	combout => \Mux72~14_combout\);

-- Location: MLABCELL_X65_Y5_N48
\Mux72~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux72~1_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux72~14_combout\)))) # (\R.curInst\(17) & ((!\Mux72~14_combout\ & ((\RegFile[12][18]~q\))) # (\Mux72~14_combout\ & (\RegFile[13][18]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux72~14_combout\)))) # (\R.curInst\(17) & ((!\Mux72~14_combout\ & ((\RegFile[14][18]~q\))) # (\Mux72~14_combout\ & (\RegFile[15][18]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][18]~q\,
	datab => \ALT_INV_RegFile[13][18]~q\,
	datac => \ALT_INV_RegFile[14][18]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux72~14_combout\,
	datag => \ALT_INV_RegFile[12][18]~q\,
	combout => \Mux72~1_combout\);

-- Location: LABCELL_X68_Y4_N24
\Mux72~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux72~13_combout\ = ( \Mux72~9_combout\ & ( \Mux72~1_combout\ & ( ((!\R.curInst\(19) & ((\Mux72~26_combout\))) # (\R.curInst\(19) & (\Mux72~5_combout\))) # (\R.curInst\(18)) ) ) ) # ( !\Mux72~9_combout\ & ( \Mux72~1_combout\ & ( (!\R.curInst\(18) & 
-- ((!\R.curInst\(19) & ((\Mux72~26_combout\))) # (\R.curInst\(19) & (\Mux72~5_combout\)))) # (\R.curInst\(18) & (((!\R.curInst\(19))))) ) ) ) # ( \Mux72~9_combout\ & ( !\Mux72~1_combout\ & ( (!\R.curInst\(18) & ((!\R.curInst\(19) & ((\Mux72~26_combout\))) # 
-- (\R.curInst\(19) & (\Mux72~5_combout\)))) # (\R.curInst\(18) & (((\R.curInst\(19))))) ) ) ) # ( !\Mux72~9_combout\ & ( !\Mux72~1_combout\ & ( (!\R.curInst\(18) & ((!\R.curInst\(19) & ((\Mux72~26_combout\))) # (\R.curInst\(19) & (\Mux72~5_combout\)))) ) ) 
-- )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001010100010000001111010011101010010111100100101011111110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(18),
	datab => \ALT_INV_Mux72~5_combout\,
	datac => \ALT_INV_R.curInst\(19),
	datad => \ALT_INV_Mux72~26_combout\,
	datae => \ALT_INV_Mux72~9_combout\,
	dataf => \ALT_INV_Mux72~1_combout\,
	combout => \Mux72~13_combout\);

-- Location: LABCELL_X74_Y6_N9
\Mux236~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux236~0_combout\ = ( \Mux72~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC\(18)))) ) ) # ( !\Mux72~13_combout\ & ( (!\vAluSrc1~1_combout\ & (\vAluSrc1~2_combout\ & \R.curPC\(18))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000001010000000000000101010100000101010101010000010101010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluSrc1~1_combout\,
	datac => \ALT_INV_vAluSrc1~2_combout\,
	datad => \ALT_INV_R.curPC\(18),
	dataf => \ALT_INV_Mux72~13_combout\,
	combout => \Mux236~0_combout\);

-- Location: FF_X74_Y6_N46
\R.aluData1[18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux236~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData1\(18));

-- Location: MLABCELL_X84_Y6_N0
\Selector14~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector14~1_combout\ = ( \R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( \R.aluData2\(18) & ( (!\R.aluOp.ALUOpXor~DUPLICATE_q\ & (!\R.aluOp.ALUOpOr~q\ & !\R.aluData1\(18))) ) ) ) # ( !\R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( \R.aluData2\(18) & ( (!\R.aluOp.ALUOpOr~q\ & 
-- ((!\R.aluOp.ALUOpXor~DUPLICATE_q\) # (\R.aluData1\(18)))) ) ) ) # ( \R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( !\R.aluData2\(18) & ( (!\R.aluData1\(18)) # ((!\R.aluOp.ALUOpXor~DUPLICATE_q\ & !\R.aluOp.ALUOpOr~q\)) ) ) ) # ( !\R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( 
-- !\R.aluData2\(18) & ( (!\R.aluData1\(18)) # ((!\R.aluOp.ALUOpXor~DUPLICATE_q\ & !\R.aluOp.ALUOpOr~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111100011111000111110001111100010001100100011001000000010000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpXor~DUPLICATE_q\,
	datab => \ALT_INV_R.aluOp.ALUOpOr~q\,
	datac => \ALT_INV_R.aluData1\(18),
	datae => \ALT_INV_R.aluOp.ALUOpAnd~DUPLICATE_q\,
	dataf => \ALT_INV_R.aluData2\(18),
	combout => \Selector14~1_combout\);

-- Location: LABCELL_X79_Y3_N9
\Selector14~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector14~2_combout\ = ( \ShiftLeft0~2_OTERM221\ & ( (!\Selector17~0_OTERM391\ & (\Selector14~1_combout\ & !\Selector16~0_OTERM393\)) ) ) # ( !\ShiftLeft0~2_OTERM221\ & ( (!\Selector17~0_OTERM391\ & \Selector14~1_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101000001010000010100000101000001010000000000000101000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector17~0_OTERM391\,
	datac => \ALT_INV_Selector14~1_combout\,
	datad => \ALT_INV_Selector16~0_OTERM393\,
	dataf => \ALT_INV_ShiftLeft0~2_OTERM221\,
	combout => \Selector14~2_combout\);

-- Location: LABCELL_X79_Y3_N42
\Selector14~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector14~3_combout\ = ( \Add2~73_sumout\ & ( (!\R.aluOp.ALUOpSub~q\ & (\Selector14~2_combout\ & ((!\R.aluOp.ALUOpAdd~q\) # (!\Add1~73_sumout\)))) ) ) # ( !\Add2~73_sumout\ & ( (\Selector14~2_combout\ & ((!\R.aluOp.ALUOpAdd~q\) # (!\Add1~73_sumout\))) ) 
-- )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110000001100110011000000100010001000000010001000100000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datab => \ALT_INV_Selector14~2_combout\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_Add1~73_sumout\,
	dataf => \ALT_INV_Add2~73_sumout\,
	combout => \Selector14~3_combout\);

-- Location: LABCELL_X77_Y4_N24
\Add3~73\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~73_sumout\ = SUM(( \R.curPC\(18) ) + ( (\R.curInst\(0) & (\R.curInst\(1) & \Mux136~0_combout\)) ) + ( \Add3~70\ ))
-- \Add3~74\ = CARRY(( \R.curPC\(18) ) + ( (\R.curInst\(0) & (\R.curInst\(1) & \Mux136~0_combout\)) ) + ( \Add3~70\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111101111111000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datac => \ALT_INV_Mux136~0_combout\,
	datad => \ALT_INV_R.curPC\(18),
	cin => \Add3~70\,
	sumout => \Add3~73_sumout\,
	cout => \Add3~74\);

-- Location: MLABCELL_X78_Y2_N12
\Comb:vJumpAdr[18]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[18]~0_combout\ = ( \Equal4~2_combout\ & ( \Add3~73_sumout\ & ( (!\R.aluCalc~q\ & (((\R.aluRes\(18))))) # (\R.aluCalc~q\ & ((!\Selector14~3_combout\) # ((\Selector14~4_combout\)))) ) ) ) # ( !\Equal4~2_combout\ & ( \Add3~73_sumout\ ) ) # ( 
-- \Equal4~2_combout\ & ( !\Add3~73_sumout\ & ( (!\R.aluCalc~q\ & (((\R.aluRes\(18))))) # (\R.aluCalc~q\ & ((!\Selector14~3_combout\) # ((\Selector14~4_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011111011101111111111111111110000111110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector14~3_combout\,
	datab => \ALT_INV_Selector14~4_combout\,
	datac => \ALT_INV_R.aluRes\(18),
	datad => \ALT_INV_R.aluCalc~q\,
	datae => \ALT_INV_Equal4~2_combout\,
	dataf => \ALT_INV_Add3~73_sumout\,
	combout => \Comb:vJumpAdr[18]~0_combout\);

-- Location: FF_X78_Y2_N13
\R.curPC[18]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[18]~0_combout\,
	asdata => \Add0~65_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(18));

-- Location: LABCELL_X81_Y6_N51
\Add0~69\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~69_sumout\ = SUM(( \R.curPC\(19) ) + ( GND ) + ( \Add0~66\ ))
-- \Add0~70\ = CARRY(( \R.curPC\(19) ) + ( GND ) + ( \Add0~66\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \ALT_INV_R.curPC\(19),
	cin => \Add0~66\,
	sumout => \Add0~69_sumout\,
	cout => \Add0~70\);

-- Location: LABCELL_X83_Y4_N24
\R.regWriteData[19]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.regWriteData[19]~feeder_combout\ = ( \Add0~69_sumout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_Add0~69_sumout\,
	combout => \R.regWriteData[19]~feeder_combout\);

-- Location: IOIBUF_X58_Y0_N75
\avm_d_readdata[11]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(11),
	o => \avm_d_readdata[11]~input_o\);

-- Location: LABCELL_X79_Y1_N48
\Comb:vRegWriteData[19]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[19]~0_combout\ = ( !\R.curInst\(13) & ( \R.curInst\(12) & ( (\avm_d_readdata[23]~input_o\ & \Comb:vRegWriteData[24]~1_combout\) ) ) ) # ( \R.curInst\(13) & ( !\R.curInst\(12) & ( (\Comb:vRegWriteData[24]~1_combout\ & 
-- \avm_d_readdata[11]~input_o\) ) ) ) # ( !\R.curInst\(13) & ( !\R.curInst\(12) & ( (\avm_d_readdata[31]~input_o\ & \Comb:vRegWriteData[24]~1_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000000000111100000101000001010000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_avm_d_readdata[23]~input_o\,
	datab => \ALT_INV_avm_d_readdata[31]~input_o\,
	datac => \ALT_INV_Comb:vRegWriteData[24]~1_combout\,
	datad => \ALT_INV_avm_d_readdata[11]~input_o\,
	datae => \ALT_INV_R.curInst\(13),
	dataf => \ALT_INV_R.curInst\(12),
	combout => \Comb:vRegWriteData[19]~0_combout\);

-- Location: LABCELL_X83_Y4_N36
\Comb:vRegWriteData[19]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[19]~1_combout\ = ( \R.memToReg~q\ & ( \Comb:vRegWriteData[19]~0_combout\ ) ) # ( !\R.memToReg~q\ & ( \Comb:vRegWriteData[19]~0_combout\ ) ) # ( !\R.memToReg~q\ & ( !\Comb:vRegWriteData[19]~0_combout\ & ( (!\R.aluCalc~q\ & 
-- (((\R.aluRes\(19))))) # (\R.aluCalc~q\ & (((!\Selector13~1_combout\)) # (\Selector13~2_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001111110101000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector13~2_combout\,
	datab => \ALT_INV_R.aluRes\(19),
	datac => \ALT_INV_Selector13~1_combout\,
	datad => \ALT_INV_R.aluCalc~q\,
	datae => \ALT_INV_R.memToReg~q\,
	dataf => \ALT_INV_Comb:vRegWriteData[19]~0_combout\,
	combout => \Comb:vRegWriteData[19]~1_combout\);

-- Location: FF_X83_Y4_N26
\R.regWriteData[19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \R.regWriteData[19]~feeder_combout\,
	asdata => \Comb:vRegWriteData[19]~1_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(19));

-- Location: FF_X73_Y3_N56
\RegFile[3][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(19),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][19]~q\);

-- Location: LABCELL_X73_Y3_N48
\Mux71~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux71~0_combout\ = ( \RegFile[7][19]~q\ & ( \R.curInst\(15) & ( (\RegFile[5][19]~q\) # (\R.curInst\(16)) ) ) ) # ( !\RegFile[7][19]~q\ & ( \R.curInst\(15) & ( (!\R.curInst\(16) & \RegFile[5][19]~q\) ) ) ) # ( \RegFile[7][19]~q\ & ( !\R.curInst\(15) & ( 
-- (!\R.curInst\(16) & (\RegFile[4][19]~q\)) # (\R.curInst\(16) & ((\RegFile[6][19]~q\))) ) ) ) # ( !\RegFile[7][19]~q\ & ( !\R.curInst\(15) & ( (!\R.curInst\(16) & (\RegFile[4][19]~q\)) # (\R.curInst\(16) & ((\RegFile[6][19]~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100010001110111010001000111011100001100000011000011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[4][19]~q\,
	datab => \ALT_INV_R.curInst\(16),
	datac => \ALT_INV_RegFile[5][19]~q\,
	datad => \ALT_INV_RegFile[6][19]~q\,
	datae => \ALT_INV_RegFile[7][19]~q\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux71~0_combout\);

-- Location: FF_X72_Y3_N58
\RegFile[1][19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[1][19]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][19]~q\);

-- Location: LABCELL_X73_Y3_N54
\Mux71~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux71~26_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (\R.curInst\(15) & (\RegFile[1][19]~q\))) # (\R.curInst\(17) & (((\Mux71~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & ((!\R.curInst\(15) & (((\RegFile[2][19]~q\)))) # 
-- (\R.curInst\(15) & (\RegFile[3][19]~q\)))) # (\R.curInst\(17) & ((((\Mux71~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000000000111010000000000000011111111110001110111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][19]~q\,
	datab => \ALT_INV_R.curInst\(15),
	datac => \ALT_INV_RegFile[2][19]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux71~0_combout\,
	datag => \ALT_INV_RegFile[1][19]~q\,
	combout => \Mux71~26_combout\);

-- Location: MLABCELL_X65_Y3_N18
\Mux71~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux71~22_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[24][19]~q\))) # (\R.curInst\(15) & (\RegFile[25][19]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[26][19]~q\))) # (\R.curInst\(15) & (\RegFile[27][19]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[27][19]~q\,
	datab => \ALT_INV_RegFile[25][19]~q\,
	datac => \ALT_INV_RegFile[26][19]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][19]~q\,
	combout => \Mux71~22_combout\);

-- Location: LABCELL_X66_Y3_N12
\Mux71~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux71~9_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux71~22_combout\))))) # (\R.curInst\(17) & (((!\Mux71~22_combout\ & (\RegFile[28][19]~q\)) # (\Mux71~22_combout\ & ((\RegFile[29][19]~q\)))))) ) ) # ( \R.curInst\(16) & ( 
-- (!\R.curInst\(17) & ((((\Mux71~22_combout\))))) # (\R.curInst\(17) & (((!\Mux71~22_combout\ & ((\RegFile[30][19]~q\))) # (\Mux71~22_combout\ & (\RegFile[31][19]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110101010111111111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[31][19]~q\,
	datac => \ALT_INV_RegFile[30][19]~q\,
	datad => \ALT_INV_RegFile[29][19]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux71~22_combout\,
	datag => \ALT_INV_RegFile[28][19]~q\,
	combout => \Mux71~9_combout\);

-- Location: LABCELL_X63_Y1_N18
\Mux71~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux71~14_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[8][19]~q\))) # (\R.curInst\(15) & (\RegFile[9][19]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[10][19]~q\))) # (\R.curInst\(15) & (\RegFile[11][19]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][19]~q\,
	datab => \ALT_INV_RegFile[11][19]~q\,
	datac => \ALT_INV_RegFile[10][19]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][19]~q\,
	combout => \Mux71~14_combout\);

-- Location: LABCELL_X63_Y3_N54
\Mux71~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux71~1_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux71~14_combout\)))) # (\R.curInst\(17) & ((!\Mux71~14_combout\ & ((\RegFile[12][19]~q\))) # (\Mux71~14_combout\ & (\RegFile[13][19]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux71~14_combout\)))) # (\R.curInst\(17) & ((!\Mux71~14_combout\ & ((\RegFile[14][19]~q\))) # (\Mux71~14_combout\ & (\RegFile[15][19]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][19]~q\,
	datab => \ALT_INV_RegFile[13][19]~q\,
	datac => \ALT_INV_RegFile[14][19]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux71~14_combout\,
	datag => \ALT_INV_RegFile[12][19]~q\,
	combout => \Mux71~1_combout\);

-- Location: MLABCELL_X72_Y1_N48
\Mux71~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux71~18_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[16][19]~q\))) # (\R.curInst\(15) & (\RegFile[17][19]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[18][19]~q\))) # (\R.curInst\(15) & (\RegFile[19][19]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[19][19]~q\,
	datab => \ALT_INV_RegFile[17][19]~q\,
	datac => \ALT_INV_RegFile[18][19]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][19]~q\,
	combout => \Mux71~18_combout\);

-- Location: MLABCELL_X72_Y1_N36
\Mux71~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux71~5_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux71~18_combout\)))) # (\R.curInst\(17) & ((!\Mux71~18_combout\ & ((\RegFile[20][19]~q\))) # (\Mux71~18_combout\ & (\RegFile[21][19]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux71~18_combout\)))) # (\R.curInst\(17) & ((!\Mux71~18_combout\ & ((\RegFile[22][19]~q\))) # (\Mux71~18_combout\ & (\RegFile[23][19]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[23][19]~q\,
	datab => \ALT_INV_RegFile[21][19]~q\,
	datac => \ALT_INV_RegFile[22][19]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux71~18_combout\,
	datag => \ALT_INV_RegFile[20][19]~q\,
	combout => \Mux71~5_combout\);

-- Location: LABCELL_X73_Y3_N39
\Mux71~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux71~13_combout\ = ( \Mux71~1_combout\ & ( \Mux71~5_combout\ & ( (!\R.curInst\(18) & (((\R.curInst\(19))) # (\Mux71~26_combout\))) # (\R.curInst\(18) & (((!\R.curInst\(19)) # (\Mux71~9_combout\)))) ) ) ) # ( !\Mux71~1_combout\ & ( \Mux71~5_combout\ & ( 
-- (!\R.curInst\(18) & (((\R.curInst\(19))) # (\Mux71~26_combout\))) # (\R.curInst\(18) & (((\Mux71~9_combout\ & \R.curInst\(19))))) ) ) ) # ( \Mux71~1_combout\ & ( !\Mux71~5_combout\ & ( (!\R.curInst\(18) & (\Mux71~26_combout\ & ((!\R.curInst\(19))))) # 
-- (\R.curInst\(18) & (((!\R.curInst\(19)) # (\Mux71~9_combout\)))) ) ) ) # ( !\Mux71~1_combout\ & ( !\Mux71~5_combout\ & ( (!\R.curInst\(18) & (\Mux71~26_combout\ & ((!\R.curInst\(19))))) # (\R.curInst\(18) & (((\Mux71~9_combout\ & \R.curInst\(19))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100010000000011011101110000001101000100110011110111011111001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux71~26_combout\,
	datab => \ALT_INV_R.curInst\(18),
	datac => \ALT_INV_Mux71~9_combout\,
	datad => \ALT_INV_R.curInst\(19),
	datae => \ALT_INV_Mux71~1_combout\,
	dataf => \ALT_INV_Mux71~5_combout\,
	combout => \Mux71~13_combout\);

-- Location: LABCELL_X74_Y6_N15
\Mux235~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux235~0_combout\ = ( \Mux71~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC\(19)))) ) ) # ( !\Mux71~13_combout\ & ( (!\vAluSrc1~1_combout\ & (\vAluSrc1~2_combout\ & \R.curPC\(19))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001000000010000000100000001010001010100010101000101010001010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluSrc1~1_combout\,
	datab => \ALT_INV_vAluSrc1~2_combout\,
	datac => \ALT_INV_R.curPC\(19),
	dataf => \ALT_INV_Mux71~13_combout\,
	combout => \Mux235~0_combout\);

-- Location: FF_X74_Y6_N41
\R.aluData1[19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux235~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData1\(19));

-- Location: IOIBUF_X36_Y0_N52
\avm_d_readdata[12]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(12),
	o => \avm_d_readdata[12]~input_o\);

-- Location: LABCELL_X79_Y8_N36
\Comb:vRegWriteData[20]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[20]~1_combout\ = ( \R.memToReg~q\ & ( \Add1~81_sumout\ & ( (!\R.curInst\(14) & ((!\R.curInst\(13)) # (\avm_d_readdata[12]~input_o\))) ) ) ) # ( !\R.memToReg~q\ & ( \Add1~81_sumout\ & ( \R.aluOp.ALUOpAdd~q\ ) ) ) # ( \R.memToReg~q\ & ( 
-- !\Add1~81_sumout\ & ( (!\R.curInst\(14) & ((!\R.curInst\(13)) # (\avm_d_readdata[12]~input_o\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100000011000001010101010101011111000000110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datab => \ALT_INV_avm_d_readdata[12]~input_o\,
	datac => \ALT_INV_R.curInst\(14),
	datad => \ALT_INV_R.curInst\(13),
	datae => \ALT_INV_R.memToReg~q\,
	dataf => \ALT_INV_Add1~81_sumout\,
	combout => \Comb:vRegWriteData[20]~1_combout\);

-- Location: LABCELL_X79_Y2_N3
\Comb:vRegWriteData[20]~2_RESYN1110\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[20]~2_RESYN1110_BDD1111\ = ( \R.curInst\(12) & ( !\avm_d_readdata[23]~input_o\ ) ) # ( !\R.curInst\(12) & ( !\avm_d_readdata[31]~input_o\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111000011110000111100001111000010101010101010101010101010101010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_avm_d_readdata[23]~input_o\,
	datac => \ALT_INV_avm_d_readdata[31]~input_o\,
	dataf => \ALT_INV_R.curInst\(12),
	combout => \Comb:vRegWriteData[20]~2_RESYN1110_BDD1111\);

-- Location: LABCELL_X79_Y2_N24
\Comb:vRegWriteData[20]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[20]~2_combout\ = ( \Comb:vRegWriteData[20]~2_RESYN1110_BDD1111\ & ( \R.curInst\(12) & ( \R.memToReg~q\ ) ) ) # ( !\Comb:vRegWriteData[20]~2_RESYN1110_BDD1111\ & ( \R.curInst\(12) & ( (\R.memToReg~q\ & ((\R.curInst\(13)) # 
-- (\R.curInst\(14)))) ) ) ) # ( \Comb:vRegWriteData[20]~2_RESYN1110_BDD1111\ & ( !\R.curInst\(12) & ( (\R.memToReg~q\ & (((!\avm_d_readdata[12]~input_o\) # (!\R.curInst\(13))) # (\R.curInst\(14)))) ) ) ) # ( !\Comb:vRegWriteData[20]~2_RESYN1110_BDD1111\ & ( 
-- !\R.curInst\(12) & ( (\R.memToReg~q\ & (((!\avm_d_readdata[12]~input_o\ & \R.curInst\(13))) # (\R.curInst\(14)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100110001001100110011000100010001001100110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(14),
	datab => \ALT_INV_R.memToReg~q\,
	datac => \ALT_INV_avm_d_readdata[12]~input_o\,
	datad => \ALT_INV_R.curInst\(13),
	datae => \ALT_INV_Comb:vRegWriteData[20]~2_RESYN1110_BDD1111\,
	dataf => \ALT_INV_R.curInst\(12),
	combout => \Comb:vRegWriteData[20]~2_combout\);

-- Location: LABCELL_X79_Y8_N48
\Comb:vRegWriteData[20]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[20]~0_combout\ = ( \Comb:vRegWriteData[20]~1_combout\ & ( !\Comb:vRegWriteData[20]~2_combout\ & ( (!\Comb:vRegWriteData[20]~3_combout\) # (\R.aluCalc~q\) ) ) ) # ( !\Comb:vRegWriteData[20]~1_combout\ & ( 
-- !\Comb:vRegWriteData[20]~2_combout\ & ( (!\Comb:vRegWriteData[20]~3_combout\) # ((\R.aluOp.ALUOpSub~q\ & (\R.aluCalc~q\ & \Add2~81_sumout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111000011110001111100111111001100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_Comb:vRegWriteData[20]~3_combout\,
	datad => \ALT_INV_Add2~81_sumout\,
	datae => \ALT_INV_Comb:vRegWriteData[20]~1_combout\,
	dataf => \ALT_INV_Comb:vRegWriteData[20]~2_combout\,
	combout => \Comb:vRegWriteData[20]~0_combout\);

-- Location: FF_X79_Y8_N14
\R.regWriteData[20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \R.regWriteData[20]~feeder_combout\,
	asdata => \Comb:vRegWriteData[20]~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(20));

-- Location: FF_X67_Y5_N31
\RegFile[6][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(20),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][20]~q\);

-- Location: FF_X68_Y3_N32
\RegFile[7][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(20),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][20]~q\);

-- Location: FF_X67_Y5_N49
\RegFile[4][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(20),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][20]~q\);

-- Location: LABCELL_X67_Y6_N6
\RegFile[5][20]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[5][20]~feeder_combout\ = ( \R.regWriteData\(20) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(20),
	combout => \RegFile[5][20]~feeder_combout\);

-- Location: FF_X67_Y6_N7
\RegFile[5][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[5][20]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][20]~q\);

-- Location: LABCELL_X68_Y3_N6
\Mux102~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux102~0_combout\ = ( \R.curInst\(21) & ( \R.curInst\(20) & ( \RegFile[7][20]~q\ ) ) ) # ( !\R.curInst\(21) & ( \R.curInst\(20) & ( \RegFile[5][20]~q\ ) ) ) # ( \R.curInst\(21) & ( !\R.curInst\(20) & ( \RegFile[6][20]~q\ ) ) ) # ( !\R.curInst\(21) & ( 
-- !\R.curInst\(20) & ( \RegFile[4][20]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111010101010101010100000000111111110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[6][20]~q\,
	datab => \ALT_INV_RegFile[7][20]~q\,
	datac => \ALT_INV_RegFile[4][20]~q\,
	datad => \ALT_INV_RegFile[5][20]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	combout => \Mux102~0_combout\);

-- Location: FF_X67_Y3_N14
\RegFile[3][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(20),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][20]~q\);

-- Location: FF_X72_Y3_N2
\RegFile[2][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(20),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][20]~q\);

-- Location: MLABCELL_X72_Y3_N54
\RegFile[1][20]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[1][20]~feeder_combout\ = ( \R.regWriteData\(20) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(20),
	combout => \RegFile[1][20]~feeder_combout\);

-- Location: FF_X72_Y3_N56
\RegFile[1][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[1][20]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][20]~q\);

-- Location: MLABCELL_X72_Y3_N0
\Mux102~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux102~26_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\RegFile[1][20]~q\ & \R.curInst\(20))))) # (\R.curInst\(22) & (\Mux102~0_combout\))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[2][20]~q\))) # 
-- (\R.curInst\(20) & (\RegFile[3][20]~q\))))) # (\R.curInst\(22) & (\Mux102~0_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000001010101000011110101010100001111010101010011001101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux102~0_combout\,
	datab => \ALT_INV_RegFile[3][20]~q\,
	datac => \ALT_INV_RegFile[2][20]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[1][20]~q\,
	combout => \Mux102~26_combout\);

-- Location: FF_X60_Y1_N38
\RegFile[21][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(20),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][20]~q\);

-- Location: FF_X65_Y2_N50
\RegFile[23][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(20),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][20]~q\);

-- Location: FF_X71_Y1_N26
\RegFile[22][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(20),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][20]~q\);

-- Location: FF_X60_Y1_N20
\RegFile[17][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(20),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][20]~q\);

-- Location: LABCELL_X60_Y1_N51
\RegFile[18][20]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[18][20]~feeder_combout\ = ( \R.regWriteData\(20) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(20),
	combout => \RegFile[18][20]~feeder_combout\);

-- Location: FF_X60_Y1_N53
\RegFile[18][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][20]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][20]~q\);

-- Location: FF_X65_Y2_N2
\RegFile[19][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(20),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][20]~q\);

-- Location: LABCELL_X57_Y2_N0
\RegFile[16][20]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[16][20]~feeder_combout\ = ( \R.regWriteData\(20) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(20),
	combout => \RegFile[16][20]~feeder_combout\);

-- Location: FF_X57_Y2_N1
\RegFile[16][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[16][20]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][20]~q\);

-- Location: LABCELL_X60_Y1_N18
\Mux102~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux102~18_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[16][20]~q\))) # (\R.curInst\(20) & (\RegFile[17][20]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & (\RegFile[18][20]~q\)) # (\R.curInst\(20) & ((\RegFile[19][20]~q\)))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001110111011101110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[17][20]~q\,
	datac => \ALT_INV_RegFile[18][20]~q\,
	datad => \ALT_INV_RegFile[19][20]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][20]~q\,
	combout => \Mux102~18_combout\);

-- Location: FF_X71_Y1_N31
\RegFile[20][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(20),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][20]~q\);

-- Location: LABCELL_X60_Y1_N36
\Mux102~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux102~5_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux102~18_combout\)))) # (\R.curInst\(22) & ((!\Mux102~18_combout\ & ((\RegFile[20][20]~q\))) # (\Mux102~18_combout\ & (\RegFile[21][20]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux102~18_combout\)))) # (\R.curInst\(22) & ((!\Mux102~18_combout\ & ((\RegFile[22][20]~q\))) # (\Mux102~18_combout\ & (\RegFile[23][20]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][20]~q\,
	datab => \ALT_INV_RegFile[23][20]~q\,
	datac => \ALT_INV_RegFile[22][20]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux102~18_combout\,
	datag => \ALT_INV_RegFile[20][20]~q\,
	combout => \Mux102~5_combout\);

-- Location: FF_X63_Y3_N26
\RegFile[15][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(20),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][20]~q\);

-- Location: FF_X63_Y1_N26
\RegFile[13][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(20),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][20]~q\);

-- Location: FF_X63_Y3_N49
\RegFile[14][20]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(20),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][20]~DUPLICATE_q\);

-- Location: FF_X63_Y1_N38
\RegFile[11][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(20),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][20]~q\);

-- Location: LABCELL_X61_Y1_N24
\RegFile[10][20]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[10][20]~feeder_combout\ = ( \R.regWriteData\(20) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(20),
	combout => \RegFile[10][20]~feeder_combout\);

-- Location: FF_X61_Y1_N25
\RegFile[10][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[10][20]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][20]~q\);

-- Location: FF_X63_Y1_N8
\RegFile[9][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(20),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][20]~q\);

-- Location: MLABCELL_X59_Y1_N57
\RegFile[8][20]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[8][20]~feeder_combout\ = ( \R.regWriteData\(20) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(20),
	combout => \RegFile[8][20]~feeder_combout\);

-- Location: FF_X59_Y1_N58
\RegFile[8][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[8][20]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][20]~q\);

-- Location: LABCELL_X63_Y1_N6
\Mux102~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux102~14_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & (\RegFile[8][20]~q\)) # (\R.curInst\(20) & ((\RegFile[9][20]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & ((\RegFile[10][20]~q\))) # (\R.curInst\(20) & (\RegFile[11][20]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110000110011111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[11][20]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[10][20]~q\,
	datad => \ALT_INV_RegFile[9][20]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][20]~q\,
	combout => \Mux102~14_combout\);

-- Location: FF_X62_Y2_N10
\RegFile[12][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(20),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][20]~q\);

-- Location: LABCELL_X63_Y1_N24
\Mux102~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux102~1_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux102~14_combout\)))) # (\R.curInst\(22) & ((!\Mux102~14_combout\ & ((\RegFile[12][20]~q\))) # (\Mux102~14_combout\ & (\RegFile[13][20]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux102~14_combout\)))) # (\R.curInst\(22) & ((!\Mux102~14_combout\ & ((\RegFile[14][20]~DUPLICATE_q\))) # (\Mux102~14_combout\ & (\RegFile[15][20]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][20]~q\,
	datab => \ALT_INV_RegFile[13][20]~q\,
	datac => \ALT_INV_RegFile[14][20]~DUPLICATE_q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux102~14_combout\,
	datag => \ALT_INV_RegFile[12][20]~q\,
	combout => \Mux102~1_combout\);

-- Location: FF_X66_Y3_N8
\RegFile[31][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(20),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][20]~q\);

-- Location: FF_X66_Y2_N38
\RegFile[29][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(20),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][20]~q\);

-- Location: LABCELL_X66_Y3_N42
\RegFile[30][20]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[30][20]~feeder_combout\ = \R.regWriteData\(20)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110011001100110011001100110011001100110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.regWriteData\(20),
	combout => \RegFile[30][20]~feeder_combout\);

-- Location: FF_X66_Y3_N43
\RegFile[30][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[30][20]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][20]~q\);

-- Location: FF_X66_Y2_N2
\RegFile[25][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(20),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][20]~q\);

-- Location: LABCELL_X60_Y2_N48
\RegFile[26][20]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[26][20]~feeder_combout\ = ( \R.regWriteData\(20) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(20),
	combout => \RegFile[26][20]~feeder_combout\);

-- Location: FF_X60_Y2_N49
\RegFile[26][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[26][20]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][20]~q\);

-- Location: FF_X66_Y2_N32
\RegFile[27][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(20),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][20]~q\);

-- Location: LABCELL_X57_Y2_N42
\RegFile[24][20]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[24][20]~feeder_combout\ = ( \R.regWriteData\(20) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(20),
	combout => \RegFile[24][20]~feeder_combout\);

-- Location: FF_X57_Y2_N43
\RegFile[24][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[24][20]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][20]~q\);

-- Location: LABCELL_X66_Y2_N0
\Mux102~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux102~22_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[24][20]~q\))) # (\R.curInst\(20) & (\RegFile[25][20]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & (\RegFile[26][20]~q\)) # (\R.curInst\(20) & ((\RegFile[27][20]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[25][20]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[26][20]~q\,
	datad => \ALT_INV_RegFile[27][20]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][20]~q\,
	combout => \Mux102~22_combout\);

-- Location: LABCELL_X66_Y3_N3
\RegFile[28][20]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[28][20]~feeder_combout\ = ( \R.regWriteData\(20) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(20),
	combout => \RegFile[28][20]~feeder_combout\);

-- Location: FF_X66_Y3_N5
\RegFile[28][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[28][20]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][20]~q\);

-- Location: LABCELL_X66_Y2_N36
\Mux102~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux102~9_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux102~22_combout\)))) # (\R.curInst\(22) & ((!\Mux102~22_combout\ & ((\RegFile[28][20]~q\))) # (\Mux102~22_combout\ & (\RegFile[29][20]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux102~22_combout\)))) # (\R.curInst\(22) & ((!\Mux102~22_combout\ & ((\RegFile[30][20]~q\))) # (\Mux102~22_combout\ & (\RegFile[31][20]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][20]~q\,
	datab => \ALT_INV_RegFile[29][20]~q\,
	datac => \ALT_INV_RegFile[30][20]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux102~22_combout\,
	datag => \ALT_INV_RegFile[28][20]~q\,
	combout => \Mux102~9_combout\);

-- Location: MLABCELL_X72_Y3_N33
\Mux102~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux102~13_combout\ = ( \Mux102~1_combout\ & ( \Mux102~9_combout\ & ( ((!\R.curInst\(24) & (\Mux102~26_combout\)) # (\R.curInst\(24) & ((\Mux102~5_combout\)))) # (\R.curInst\(23)) ) ) ) # ( !\Mux102~1_combout\ & ( \Mux102~9_combout\ & ( (!\R.curInst\(24) 
-- & (\Mux102~26_combout\ & ((!\R.curInst\(23))))) # (\R.curInst\(24) & (((\R.curInst\(23)) # (\Mux102~5_combout\)))) ) ) ) # ( \Mux102~1_combout\ & ( !\Mux102~9_combout\ & ( (!\R.curInst\(24) & (((\R.curInst\(23))) # (\Mux102~26_combout\))) # 
-- (\R.curInst\(24) & (((\Mux102~5_combout\ & !\R.curInst\(23))))) ) ) ) # ( !\Mux102~1_combout\ & ( !\Mux102~9_combout\ & ( (!\R.curInst\(23) & ((!\R.curInst\(24) & (\Mux102~26_combout\)) # (\R.curInst\(24) & ((\Mux102~5_combout\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100011100000000010001111100110001000111001100110100011111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux102~26_combout\,
	datab => \ALT_INV_R.curInst\(24),
	datac => \ALT_INV_Mux102~5_combout\,
	datad => \ALT_INV_R.curInst\(23),
	datae => \ALT_INV_Mux102~1_combout\,
	dataf => \ALT_INV_Mux102~9_combout\,
	combout => \Mux102~13_combout\);

-- Location: LABCELL_X73_Y5_N54
\NxR.aluData2[20]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[20]~1_combout\ = ( \vAluSrc2~1_combout\ & ( (\Mux134~0_combout\ & \Equal4~1_combout\) ) ) # ( !\vAluSrc2~1_combout\ & ( \Mux102~13_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111000000001111111100000011000000110000001100000011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Mux134~0_combout\,
	datac => \ALT_INV_Equal4~1_combout\,
	datad => \ALT_INV_Mux102~13_combout\,
	dataf => \ALT_INV_vAluSrc2~1_combout\,
	combout => \NxR.aluData2[20]~1_combout\);

-- Location: FF_X73_Y5_N40
\R.aluData2[20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \NxR.aluData2[20]~1_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData2\(20));

-- Location: LABCELL_X77_Y3_N21
\Selector2~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector2~3_combout\ = ( \Add1~121_sumout\ & ( \Add2~121_sumout\ & ( ((\R.aluOp.ALUOpAdd~q\) # (\R.aluOp.ALUOpSub~q\)) # (\Selector2~2_combout\) ) ) ) # ( !\Add1~121_sumout\ & ( \Add2~121_sumout\ & ( (\R.aluOp.ALUOpSub~q\) # (\Selector2~2_combout\) ) ) ) 
-- # ( \Add1~121_sumout\ & ( !\Add2~121_sumout\ & ( (\R.aluOp.ALUOpAdd~q\) # (\Selector2~2_combout\) ) ) ) # ( !\Add1~121_sumout\ & ( !\Add2~121_sumout\ & ( \Selector2~2_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101010101011111111101011111010111110101111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector2~2_combout\,
	datac => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datad => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datae => \ALT_INV_Add1~121_sumout\,
	dataf => \ALT_INV_Add2~121_sumout\,
	combout => \Selector2~3_combout\);

-- Location: FF_X77_Y3_N22
\R.aluRes[30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector2~3_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(30));

-- Location: IOIBUF_X54_Y0_N52
\avm_d_readdata[6]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(6),
	o => \avm_d_readdata[6]~input_o\);

-- Location: LABCELL_X79_Y1_N54
\Comb:vRegWriteData[30]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[30]~1_combout\ = ( !\R.curInst\(13) & ( \R.curInst\(12) & ( (!\R.curInst\(14) & \avm_d_readdata[23]~input_o\) ) ) ) # ( \R.curInst\(13) & ( !\R.curInst\(12) & ( (!\R.curInst\(14) & \avm_d_readdata[6]~input_o\) ) ) ) # ( 
-- !\R.curInst\(13) & ( !\R.curInst\(12) & ( (!\R.curInst\(14) & \avm_d_readdata[31]~input_o\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000010101010001000100010001000001010000010100000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(14),
	datab => \ALT_INV_avm_d_readdata[6]~input_o\,
	datac => \ALT_INV_avm_d_readdata[23]~input_o\,
	datad => \ALT_INV_avm_d_readdata[31]~input_o\,
	datae => \ALT_INV_R.curInst\(13),
	dataf => \ALT_INV_R.curInst\(12),
	combout => \Comb:vRegWriteData[30]~1_combout\);

-- Location: MLABCELL_X78_Y5_N51
\Comb:vRegWriteData[30]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[30]~2_combout\ = ( \Comb:vRegWriteData[30]~1_combout\ & ( (!\R.memToReg~q\ & (!\Selector2~2_combout\ & ((!\R.aluOp.ALUOpAdd~q\) # (!\Add1~121_sumout\)))) ) ) # ( !\Comb:vRegWriteData[30]~1_combout\ & ( ((!\Selector2~2_combout\ & 
-- ((!\R.aluOp.ALUOpAdd~q\) # (!\Add1~121_sumout\)))) # (\R.memToReg~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111110101010101111111010101010110101000000000001010100000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.memToReg~q\,
	datab => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datac => \ALT_INV_Add1~121_sumout\,
	datad => \ALT_INV_Selector2~2_combout\,
	dataf => \ALT_INV_Comb:vRegWriteData[30]~1_combout\,
	combout => \Comb:vRegWriteData[30]~2_combout\);

-- Location: LABCELL_X80_Y5_N48
\Comb:vRegWriteData[30]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[30]~0_combout\ = ( \Comb:vRegWriteData[30]~2_combout\ & ( \Add2~121_sumout\ & ( (!\R.memToReg~q\ & ((!\R.aluCalc~q\ & ((\R.aluRes\(30)))) # (\R.aluCalc~q\ & (\R.aluOp.ALUOpSub~q\)))) ) ) ) # ( !\Comb:vRegWriteData[30]~2_combout\ & ( 
-- \Add2~121_sumout\ & ( ((\R.aluRes\(30)) # (\R.aluCalc~q\)) # (\R.memToReg~q\) ) ) ) # ( \Comb:vRegWriteData[30]~2_combout\ & ( !\Add2~121_sumout\ & ( (!\R.memToReg~q\ & (!\R.aluCalc~q\ & \R.aluRes\(30))) ) ) ) # ( !\Comb:vRegWriteData[30]~2_combout\ & ( 
-- !\Add2~121_sumout\ & ( ((\R.aluRes\(30)) # (\R.aluCalc~q\)) # (\R.memToReg~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011111111111111000000001100000000111111111111110000010011000100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datab => \ALT_INV_R.memToReg~q\,
	datac => \ALT_INV_R.aluCalc~q\,
	datad => \ALT_INV_R.aluRes\(30),
	datae => \ALT_INV_Comb:vRegWriteData[30]~2_combout\,
	dataf => \ALT_INV_Add2~121_sumout\,
	combout => \Comb:vRegWriteData[30]~0_combout\);

-- Location: FF_X81_Y5_N56
\R.regWriteData[30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Add0~113_sumout\,
	asdata => \Comb:vRegWriteData[30]~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(30));

-- Location: FF_X64_Y2_N26
\RegFile[23][30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(30),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][30]~q\);

-- Location: LABCELL_X64_Y2_N48
\Mux60~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux60~18_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & (\RegFile[16][30]~q\)) # (\R.curInst\(15) & ((\RegFile[17][30]~q\)))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & ((\RegFile[18][30]~q\))) # (\R.curInst\(15) & (\RegFile[19][30]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001010101111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[19][30]~q\,
	datac => \ALT_INV_RegFile[18][30]~q\,
	datad => \ALT_INV_RegFile[17][30]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][30]~q\,
	combout => \Mux60~18_combout\);

-- Location: LABCELL_X64_Y2_N24
\Mux60~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux60~5_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux60~18_combout\)))) # (\R.curInst\(17) & ((!\Mux60~18_combout\ & ((\RegFile[20][30]~q\))) # (\Mux60~18_combout\ & (\RegFile[21][30]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux60~18_combout\)))) # (\R.curInst\(17) & ((!\Mux60~18_combout\ & ((\RegFile[22][30]~q\))) # (\Mux60~18_combout\ & (\RegFile[23][30]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[23][30]~q\,
	datab => \ALT_INV_RegFile[21][30]~q\,
	datac => \ALT_INV_RegFile[22][30]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux60~18_combout\,
	datag => \ALT_INV_RegFile[20][30]~q\,
	combout => \Mux60~5_combout\);

-- Location: FF_X66_Y3_N56
\RegFile[30][30]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[30][30]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][30]~DUPLICATE_q\);

-- Location: LABCELL_X66_Y2_N6
\Mux60~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux60~22_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[24][30]~q\))) # (\R.curInst\(15) & (\RegFile[25][30]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[26][30]~q\))) # (\R.curInst\(15) & (\RegFile[27][30]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[27][30]~q\,
	datab => \ALT_INV_RegFile[25][30]~q\,
	datac => \ALT_INV_RegFile[26][30]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][30]~q\,
	combout => \Mux60~22_combout\);

-- Location: LABCELL_X66_Y3_N30
\Mux60~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux60~9_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux60~22_combout\))))) # (\R.curInst\(17) & (((!\Mux60~22_combout\ & (\RegFile[28][30]~q\)) # (\Mux60~22_combout\ & ((\RegFile[29][30]~q\)))))) ) ) # ( \R.curInst\(16) & ( 
-- (!\R.curInst\(17) & ((((\Mux60~22_combout\))))) # (\R.curInst\(17) & (((!\Mux60~22_combout\ & ((\RegFile[30][30]~DUPLICATE_q\))) # (\Mux60~22_combout\ & (\RegFile[31][30]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110101010111111111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[31][30]~q\,
	datac => \ALT_INV_RegFile[30][30]~DUPLICATE_q\,
	datad => \ALT_INV_RegFile[29][30]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux60~22_combout\,
	datag => \ALT_INV_RegFile[28][30]~q\,
	combout => \Mux60~9_combout\);

-- Location: LABCELL_X67_Y3_N54
\Mux60~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux60~0_combout\ = ( \RegFile[7][30]~q\ & ( \R.curInst\(15) & ( (\R.curInst\(16)) # (\RegFile[5][30]~q\) ) ) ) # ( !\RegFile[7][30]~q\ & ( \R.curInst\(15) & ( (\RegFile[5][30]~q\ & !\R.curInst\(16)) ) ) ) # ( \RegFile[7][30]~q\ & ( !\R.curInst\(15) & ( 
-- (!\R.curInst\(16) & (\RegFile[4][30]~q\)) # (\R.curInst\(16) & ((\RegFile[6][30]~q\))) ) ) ) # ( !\RegFile[7][30]~q\ & ( !\R.curInst\(15) & ( (!\R.curInst\(16) & (\RegFile[4][30]~q\)) # (\R.curInst\(16) & ((\RegFile[6][30]~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010100001111010101010000111100110011000000000011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[4][30]~q\,
	datab => \ALT_INV_RegFile[5][30]~q\,
	datac => \ALT_INV_RegFile[6][30]~q\,
	datad => \ALT_INV_R.curInst\(16),
	datae => \ALT_INV_RegFile[7][30]~q\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux60~0_combout\);

-- Location: LABCELL_X67_Y3_N36
\Mux60~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux60~26_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((\RegFile[1][30]~q\ & ((\R.curInst\(15))))))) # (\R.curInst\(17) & (\Mux60~0_combout\)) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & (\RegFile[2][30]~q\)) # 
-- (\R.curInst\(15) & ((\RegFile[3][30]~q\)))))) # (\R.curInst\(17) & (\Mux60~0_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0001000100010001000111010001110100011101000111010001000111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux60~0_combout\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[2][30]~q\,
	datad => \ALT_INV_RegFile[3][30]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[1][30]~q\,
	combout => \Mux60~26_combout\);

-- Location: LABCELL_X70_Y2_N12
\Mux60~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux60~14_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & (\RegFile[8][30]~q\)) # (\R.curInst\(15) & ((\RegFile[9][30]~q\))))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & ((\RegFile[10][30]~q\))) # (\R.curInst\(15) & (\RegFile[11][30]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110000110011111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[11][30]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[10][30]~q\,
	datad => \ALT_INV_RegFile[9][30]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][30]~q\,
	combout => \Mux60~14_combout\);

-- Location: LABCELL_X70_Y2_N54
\Mux60~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux60~1_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux60~14_combout\)))) # (\R.curInst\(17) & ((!\Mux60~14_combout\ & ((\RegFile[12][30]~q\))) # (\Mux60~14_combout\ & (\RegFile[13][30]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux60~14_combout\)))) # (\R.curInst\(17) & ((!\Mux60~14_combout\ & ((\RegFile[14][30]~q\))) # (\Mux60~14_combout\ & (\RegFile[15][30]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][30]~q\,
	datab => \ALT_INV_RegFile[13][30]~q\,
	datac => \ALT_INV_RegFile[14][30]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux60~14_combout\,
	datag => \ALT_INV_RegFile[12][30]~q\,
	combout => \Mux60~1_combout\);

-- Location: LABCELL_X67_Y3_N24
\Mux60~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux60~13_combout\ = ( \Mux60~26_combout\ & ( \Mux60~1_combout\ & ( (!\R.curInst\(19)) # ((!\R.curInst\(18) & (\Mux60~5_combout\)) # (\R.curInst\(18) & ((\Mux60~9_combout\)))) ) ) ) # ( !\Mux60~26_combout\ & ( \Mux60~1_combout\ & ( (!\R.curInst\(18) & 
-- (\Mux60~5_combout\ & ((\R.curInst\(19))))) # (\R.curInst\(18) & (((!\R.curInst\(19)) # (\Mux60~9_combout\)))) ) ) ) # ( \Mux60~26_combout\ & ( !\Mux60~1_combout\ & ( (!\R.curInst\(18) & (((!\R.curInst\(19))) # (\Mux60~5_combout\))) # (\R.curInst\(18) & 
-- (((\Mux60~9_combout\ & \R.curInst\(19))))) ) ) ) # ( !\Mux60~26_combout\ & ( !\Mux60~1_combout\ & ( (\R.curInst\(19) & ((!\R.curInst\(18) & (\Mux60~5_combout\)) # (\R.curInst\(18) & ((\Mux60~9_combout\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000100111101010100010011101010101001001111111111100100111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(18),
	datab => \ALT_INV_Mux60~5_combout\,
	datac => \ALT_INV_Mux60~9_combout\,
	datad => \ALT_INV_R.curInst\(19),
	datae => \ALT_INV_Mux60~26_combout\,
	dataf => \ALT_INV_Mux60~1_combout\,
	combout => \Mux60~13_combout\);

-- Location: LABCELL_X73_Y5_N30
\Mux224~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux224~0_combout\ = ( \Mux60~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC[30]~DUPLICATE_q\))) ) ) # ( !\Mux60~13_combout\ & ( (\vAluSrc1~2_combout\ & (\R.curPC[30]~DUPLICATE_q\ & !\vAluSrc1~1_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000000000001010000000010101111000000001010111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluSrc1~2_combout\,
	datac => \ALT_INV_R.curPC[30]~DUPLICATE_q\,
	datad => \ALT_INV_vAluSrc1~1_combout\,
	dataf => \ALT_INV_Mux60~13_combout\,
	combout => \Mux224~0_combout\);

-- Location: LABCELL_X73_Y5_N45
\ShiftRight0~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight0~0_combout\ = ( \NxR.aluData2[1]~17_combout\ & ( (\Mux223~0_combout\ & !\NxR.aluData2[0]~16_combout\) ) ) # ( !\NxR.aluData2[1]~17_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (\Mux225~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & 
-- ((\Mux224~0_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010100001111010101010000111100110011000000000011001100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux225~0_combout\,
	datab => \ALT_INV_Mux223~0_combout\,
	datac => \ALT_INV_Mux224~0_combout\,
	datad => \ALT_INV_NxR.aluData2[0]~16_combout\,
	dataf => \ALT_INV_NxR.aluData2[1]~17_combout\,
	combout => \ShiftRight0~0_combout\);

-- Location: FF_X73_Y5_N46
\ShiftRight0~0_NEW_REG16\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight0~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight0~0_OTERM17\);

-- Location: LABCELL_X75_Y5_N18
\Selector7~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector7~0_combout\ = ( \ShiftRight0~0_OTERM17\ & ( !\R.aluData2\(3) & ( (\R.aluOp.ALUOpSRL~q\ & ((\R.aluData2\(2)) # (\ShiftRight1~12_OTERM57\))) ) ) ) # ( !\ShiftRight0~0_OTERM17\ & ( !\R.aluData2\(3) & ( (\ShiftRight1~12_OTERM57\ & (!\R.aluData2\(2) 
-- & \R.aluOp.ALUOpSRL~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110000000000000011111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_ShiftRight1~12_OTERM57\,
	datac => \ALT_INV_R.aluData2\(2),
	datad => \ALT_INV_R.aluOp.ALUOpSRL~q\,
	datae => \ALT_INV_ShiftRight0~0_OTERM17\,
	dataf => \ALT_INV_R.aluData2\(3),
	combout => \Selector7~0_combout\);

-- Location: LABCELL_X74_Y3_N6
\ShiftLeft0~42\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~42_combout\ = ( \NxR.aluData2[0]~16_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( \Mux232~0_combout\ ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( \Mux231~0_combout\ ) ) ) # ( \NxR.aluData2[0]~16_combout\ & ( 
-- !\NxR.aluData2[1]~17_combout\ & ( \Mux230~0_combout\ ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( !\NxR.aluData2[1]~17_combout\ & ( \Mux229~0_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111010101010101010100110011001100110000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux230~0_combout\,
	datab => \ALT_INV_Mux231~0_combout\,
	datac => \ALT_INV_Mux229~0_combout\,
	datad => \ALT_INV_Mux232~0_combout\,
	datae => \ALT_INV_NxR.aluData2[0]~16_combout\,
	dataf => \ALT_INV_NxR.aluData2[1]~17_combout\,
	combout => \ShiftLeft0~42_combout\);

-- Location: FF_X74_Y3_N7
\ShiftLeft0~42_NEW_REG40\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~42_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~42_OTERM41\);

-- Location: MLABCELL_X82_Y4_N36
\ShiftLeft0~43\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~43_combout\ = ( \ShiftLeft0~42_OTERM41\ & ( \ShiftLeft0~26_OTERM739\ & ( (!\R.aluData2\(2)) # ((!\R.aluData2\(3) & (\ShiftLeft0~34_OTERM299\)) # (\R.aluData2\(3) & ((\ShiftLeft0~18_OTERM289\)))) ) ) ) # ( !\ShiftLeft0~42_OTERM41\ & ( 
-- \ShiftLeft0~26_OTERM739\ & ( (!\R.aluData2\(3) & (\ShiftLeft0~34_OTERM299\ & ((\R.aluData2\(2))))) # (\R.aluData2\(3) & (((!\R.aluData2\(2)) # (\ShiftLeft0~18_OTERM289\)))) ) ) ) # ( \ShiftLeft0~42_OTERM41\ & ( !\ShiftLeft0~26_OTERM739\ & ( 
-- (!\R.aluData2\(3) & (((!\R.aluData2\(2))) # (\ShiftLeft0~34_OTERM299\))) # (\R.aluData2\(3) & (((\ShiftLeft0~18_OTERM289\ & \R.aluData2\(2))))) ) ) ) # ( !\ShiftLeft0~42_OTERM41\ & ( !\ShiftLeft0~26_OTERM739\ & ( (\R.aluData2\(2) & ((!\R.aluData2\(3) & 
-- (\ShiftLeft0~34_OTERM299\)) # (\R.aluData2\(3) & ((\ShiftLeft0~18_OTERM289\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001000111110011000100011100110011010001111111111101000111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~34_OTERM299\,
	datab => \ALT_INV_R.aluData2\(3),
	datac => \ALT_INV_ShiftLeft0~18_OTERM289\,
	datad => \ALT_INV_R.aluData2\(2),
	datae => \ALT_INV_ShiftLeft0~42_OTERM41\,
	dataf => \ALT_INV_ShiftLeft0~26_OTERM739\,
	combout => \ShiftLeft0~43_combout\);

-- Location: MLABCELL_X82_Y5_N54
\Selector7~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector7~1_combout\ = ( \R.aluOp.ALUOpSLL~q\ & ( \ShiftLeft0~43_combout\ & ( !\R.aluData2\(4) ) ) ) # ( !\R.aluOp.ALUOpSLL~q\ & ( \ShiftLeft0~43_combout\ & ( (!\R.aluData2\(4) & (((\R.aluOp.ALUOpSRA~q\ & \ShiftRight1~55_combout\)) # 
-- (\Selector7~0_combout\))) ) ) ) # ( \R.aluOp.ALUOpSLL~q\ & ( !\ShiftLeft0~43_combout\ & ( (!\R.aluData2\(4) & (((\R.aluOp.ALUOpSRA~q\ & \ShiftRight1~55_combout\)) # (\Selector7~0_combout\))) ) ) ) # ( !\R.aluOp.ALUOpSLL~q\ & ( !\ShiftLeft0~43_combout\ & ( 
-- (!\R.aluData2\(4) & (((\R.aluOp.ALUOpSRA~q\ & \ShiftRight1~55_combout\)) # (\Selector7~0_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001010101010000000101010101000000010101010101010101010101010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(4),
	datab => \ALT_INV_R.aluOp.ALUOpSRA~q\,
	datac => \ALT_INV_ShiftRight1~55_combout\,
	datad => \ALT_INV_Selector7~0_combout\,
	datae => \ALT_INV_R.aluOp.ALUOpSLL~q\,
	dataf => \ALT_INV_ShiftLeft0~43_combout\,
	combout => \Selector7~1_combout\);

-- Location: MLABCELL_X82_Y5_N18
\Comb:vRegWriteData[25]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[25]~3_combout\ = ( \R.aluRes\(25) & ( (!\Selector7~1_combout\ & (\R.aluCalc~q\ & !\Selector7~5_combout\)) ) ) # ( !\R.aluRes\(25) & ( (!\R.aluCalc~q\ & (((!\R.memToReg~q\)))) # (\R.aluCalc~q\ & (!\Selector7~1_combout\ & 
-- ((!\Selector7~5_combout\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1100101011000000000010100000000011001010110000000000101000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector7~1_combout\,
	datab => \ALT_INV_R.memToReg~q\,
	datac => \ALT_INV_R.aluCalc~q\,
	datad => \ALT_INV_Selector7~5_combout\,
	datae => \ALT_INV_R.aluRes\(25),
	combout => \Comb:vRegWriteData[25]~3_combout\);

-- Location: IOIBUF_X88_Y0_N19
\avm_d_readdata[1]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(1),
	o => \avm_d_readdata[1]~input_o\);

-- Location: MLABCELL_X82_Y5_N12
\Comb:vRegWriteData[25]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[25]~1_combout\ = ( \avm_d_readdata[1]~input_o\ & ( \Add1~101_sumout\ & ( (!\R.memToReg~q\ & ((\R.aluOp.ALUOpAdd~q\))) # (\R.memToReg~q\ & (!\R.curInst\(14))) ) ) ) # ( !\avm_d_readdata[1]~input_o\ & ( \Add1~101_sumout\ & ( 
-- (!\R.memToReg~q\ & (((\R.aluOp.ALUOpAdd~q\)))) # (\R.memToReg~q\ & (!\R.curInst\(14) & ((!\R.curInst\(13))))) ) ) ) # ( \avm_d_readdata[1]~input_o\ & ( !\Add1~101_sumout\ & ( (!\R.curInst\(14) & \R.memToReg~q\) ) ) ) # ( !\avm_d_readdata[1]~input_o\ & ( 
-- !\Add1~101_sumout\ & ( (!\R.curInst\(14) & (!\R.curInst\(13) & \R.memToReg~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000010100000000000001010101000110011101000000011001110101010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(14),
	datab => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datac => \ALT_INV_R.curInst\(13),
	datad => \ALT_INV_R.memToReg~q\,
	datae => \ALT_INV_avm_d_readdata[1]~input_o\,
	dataf => \ALT_INV_Add1~101_sumout\,
	combout => \Comb:vRegWriteData[25]~1_combout\);

-- Location: LABCELL_X79_Y1_N9
\Comb:vRegWriteData[25]~2_RESYN1106\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[25]~2_RESYN1106_BDD1107\ = ( \R.curInst\(12) & ( !\avm_d_readdata[23]~input_o\ ) ) # ( !\R.curInst\(12) & ( !\avm_d_readdata[31]~input_o\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1100110011001100110011001100110010101010101010101010101010101010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_avm_d_readdata[23]~input_o\,
	datab => \ALT_INV_avm_d_readdata[31]~input_o\,
	dataf => \ALT_INV_R.curInst\(12),
	combout => \Comb:vRegWriteData[25]~2_RESYN1106_BDD1107\);

-- Location: LABCELL_X79_Y1_N42
\Comb:vRegWriteData[25]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[25]~2_combout\ = ( \avm_d_readdata[1]~input_o\ & ( \Comb:vRegWriteData[25]~2_RESYN1106_BDD1107\ & ( (\R.memToReg~q\ & (((!\R.curInst\(13)) # (\R.curInst\(12))) # (\R.curInst\(14)))) ) ) ) # ( !\avm_d_readdata[1]~input_o\ & ( 
-- \Comb:vRegWriteData[25]~2_RESYN1106_BDD1107\ & ( \R.memToReg~q\ ) ) ) # ( \avm_d_readdata[1]~input_o\ & ( !\Comb:vRegWriteData[25]~2_RESYN1106_BDD1107\ & ( (\R.memToReg~q\ & (((\R.curInst\(13) & \R.curInst\(12))) # (\R.curInst\(14)))) ) ) ) # ( 
-- !\avm_d_readdata[1]~input_o\ & ( !\Comb:vRegWriteData[25]~2_RESYN1106_BDD1107\ & ( (\R.memToReg~q\ & ((\R.curInst\(13)) # (\R.curInst\(14)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001110111000000000101011100000000111111110000000011011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(14),
	datab => \ALT_INV_R.curInst\(13),
	datac => \ALT_INV_R.curInst\(12),
	datad => \ALT_INV_R.memToReg~q\,
	datae => \ALT_INV_avm_d_readdata[1]~input_o\,
	dataf => \ALT_INV_Comb:vRegWriteData[25]~2_RESYN1106_BDD1107\,
	combout => \Comb:vRegWriteData[25]~2_combout\);

-- Location: MLABCELL_X82_Y5_N6
\Comb:vRegWriteData[25]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[25]~0_combout\ = ( \R.aluOp.ALUOpSub~q\ & ( !\Comb:vRegWriteData[25]~2_combout\ & ( (!\Comb:vRegWriteData[25]~3_combout\) # ((\R.aluCalc~q\ & ((\Comb:vRegWriteData[25]~1_combout\) # (\Add2~101_sumout\)))) ) ) ) # ( 
-- !\R.aluOp.ALUOpSub~q\ & ( !\Comb:vRegWriteData[25]~2_combout\ & ( (!\Comb:vRegWriteData[25]~3_combout\) # ((\R.aluCalc~q\ & \Comb:vRegWriteData[25]~1_combout\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010101010101111101010111010111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Comb:vRegWriteData[25]~3_combout\,
	datab => \ALT_INV_Add2~101_sumout\,
	datac => \ALT_INV_R.aluCalc~q\,
	datad => \ALT_INV_Comb:vRegWriteData[25]~1_combout\,
	datae => \ALT_INV_R.aluOp.ALUOpSub~q\,
	dataf => \ALT_INV_Comb:vRegWriteData[25]~2_combout\,
	combout => \Comb:vRegWriteData[25]~0_combout\);

-- Location: FF_X81_Y5_N41
\R.regWriteData[25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Add0~93_sumout\,
	asdata => \Comb:vRegWriteData[25]~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(25));

-- Location: FF_X67_Y1_N2
\RegFile[31][25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(25),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][25]~q\);

-- Location: LABCELL_X67_Y1_N48
\Mux65~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux65~22_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[24][25]~q\))) # (\R.curInst\(15) & (\RegFile[25][25]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & (\RegFile[26][25]~q\)) # (\R.curInst\(15) & ((\RegFile[27][25]~q\))))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[25][25]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[26][25]~q\,
	datad => \ALT_INV_RegFile[27][25]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][25]~q\,
	combout => \Mux65~22_combout\);

-- Location: LABCELL_X67_Y1_N0
\Mux65~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux65~9_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux65~22_combout\)))) # (\R.curInst\(17) & ((!\Mux65~22_combout\ & ((\RegFile[28][25]~q\))) # (\Mux65~22_combout\ & (\RegFile[29][25]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux65~22_combout\)))) # (\R.curInst\(17) & ((!\Mux65~22_combout\ & ((\RegFile[30][25]~q\))) # (\Mux65~22_combout\ & (\RegFile[31][25]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][25]~q\,
	datab => \ALT_INV_RegFile[29][25]~q\,
	datac => \ALT_INV_RegFile[30][25]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux65~22_combout\,
	datag => \ALT_INV_RegFile[28][25]~q\,
	combout => \Mux65~9_combout\);

-- Location: LABCELL_X64_Y2_N12
\Mux65~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux65~18_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[16][25]~q\))) # (\R.curInst\(15) & (\RegFile[17][25]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[18][25]~q\))) # (\R.curInst\(15) & (\RegFile[19][25]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[17][25]~q\,
	datab => \ALT_INV_RegFile[19][25]~q\,
	datac => \ALT_INV_RegFile[18][25]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][25]~q\,
	combout => \Mux65~18_combout\);

-- Location: LABCELL_X64_Y2_N6
\Mux65~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux65~5_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux65~18_combout\)))) # (\R.curInst\(17) & ((!\Mux65~18_combout\ & ((\RegFile[20][25]~q\))) # (\Mux65~18_combout\ & (\RegFile[21][25]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux65~18_combout\)))) # (\R.curInst\(17) & ((!\Mux65~18_combout\ & ((\RegFile[22][25]~q\))) # (\Mux65~18_combout\ & (\RegFile[23][25]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][25]~q\,
	datab => \ALT_INV_RegFile[23][25]~q\,
	datac => \ALT_INV_RegFile[22][25]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux65~18_combout\,
	datag => \ALT_INV_RegFile[20][25]~q\,
	combout => \Mux65~5_combout\);

-- Location: LABCELL_X68_Y3_N12
\Mux65~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux65~0_combout\ = ( \RegFile[7][25]~q\ & ( \R.curInst\(15) & ( (\RegFile[5][25]~q\) # (\R.curInst\(16)) ) ) ) # ( !\RegFile[7][25]~q\ & ( \R.curInst\(15) & ( (!\R.curInst\(16) & \RegFile[5][25]~q\) ) ) ) # ( \RegFile[7][25]~q\ & ( !\R.curInst\(15) & ( 
-- (!\R.curInst\(16) & (\RegFile[4][25]~q\)) # (\R.curInst\(16) & ((\RegFile[6][25]~q\))) ) ) ) # ( !\RegFile[7][25]~q\ & ( !\R.curInst\(15) & ( (!\R.curInst\(16) & (\RegFile[4][25]~q\)) # (\R.curInst\(16) & ((\RegFile[6][25]~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101001101010011010100110101001100000000111100000000111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[4][25]~q\,
	datab => \ALT_INV_RegFile[6][25]~q\,
	datac => \ALT_INV_R.curInst\(16),
	datad => \ALT_INV_RegFile[5][25]~q\,
	datae => \ALT_INV_RegFile[7][25]~q\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux65~0_combout\);

-- Location: LABCELL_X68_Y3_N0
\Mux65~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux65~26_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (\RegFile[1][25]~q\ & (\R.curInst\(15)))) # (\R.curInst\(17) & (((\Mux65~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & ((!\R.curInst\(15) & (((\RegFile[2][25]~q\)))) # 
-- (\R.curInst\(15) & (\RegFile[3][25]~q\)))) # (\R.curInst\(17) & ((((\Mux65~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001100000011000100010000110011001111110011111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][25]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[2][25]~q\,
	datad => \ALT_INV_R.curInst\(15),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux65~0_combout\,
	datag => \ALT_INV_RegFile[1][25]~q\,
	combout => \Mux65~26_combout\);

-- Location: LABCELL_X68_Y2_N36
\Mux65~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux65~14_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[8][25]~q\))) # (\R.curInst\(15) & (\RegFile[9][25]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[10][25]~q\))) # (\R.curInst\(15) & (\RegFile[11][25]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[11][25]~q\,
	datab => \ALT_INV_RegFile[9][25]~q\,
	datac => \ALT_INV_RegFile[10][25]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][25]~q\,
	combout => \Mux65~14_combout\);

-- Location: LABCELL_X68_Y2_N48
\Mux65~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux65~1_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux65~14_combout\)))) # (\R.curInst\(17) & ((!\Mux65~14_combout\ & ((\RegFile[12][25]~q\))) # (\Mux65~14_combout\ & (\RegFile[13][25]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux65~14_combout\)))) # (\R.curInst\(17) & ((!\Mux65~14_combout\ & ((\RegFile[14][25]~q\))) # (\Mux65~14_combout\ & (\RegFile[15][25]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][25]~q\,
	datab => \ALT_INV_RegFile[13][25]~q\,
	datac => \ALT_INV_RegFile[14][25]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux65~14_combout\,
	datag => \ALT_INV_RegFile[12][25]~q\,
	combout => \Mux65~1_combout\);

-- Location: LABCELL_X68_Y2_N18
\Mux65~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux65~13_combout\ = ( \Mux65~26_combout\ & ( \Mux65~1_combout\ & ( (!\R.curInst\(19)) # ((!\R.curInst\(18) & ((\Mux65~5_combout\))) # (\R.curInst\(18) & (\Mux65~9_combout\))) ) ) ) # ( !\Mux65~26_combout\ & ( \Mux65~1_combout\ & ( (!\R.curInst\(19) & 
-- (\R.curInst\(18))) # (\R.curInst\(19) & ((!\R.curInst\(18) & ((\Mux65~5_combout\))) # (\R.curInst\(18) & (\Mux65~9_combout\)))) ) ) ) # ( \Mux65~26_combout\ & ( !\Mux65~1_combout\ & ( (!\R.curInst\(19) & (!\R.curInst\(18))) # (\R.curInst\(19) & 
-- ((!\R.curInst\(18) & ((\Mux65~5_combout\))) # (\R.curInst\(18) & (\Mux65~9_combout\)))) ) ) ) # ( !\Mux65~26_combout\ & ( !\Mux65~1_combout\ & ( (\R.curInst\(19) & ((!\R.curInst\(18) & ((\Mux65~5_combout\))) # (\R.curInst\(18) & (\Mux65~9_combout\)))) ) ) 
-- )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000101000101100010011100110100100011011001111010101111101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(19),
	datab => \ALT_INV_R.curInst\(18),
	datac => \ALT_INV_Mux65~9_combout\,
	datad => \ALT_INV_Mux65~5_combout\,
	datae => \ALT_INV_Mux65~26_combout\,
	dataf => \ALT_INV_Mux65~1_combout\,
	combout => \Mux65~13_combout\);

-- Location: LABCELL_X74_Y3_N51
\Mux229~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux229~0_combout\ = ( \Mux65~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC\(25)))) ) ) # ( !\Mux65~13_combout\ & ( (\vAluSrc1~2_combout\ & (\R.curPC\(25) & !\vAluSrc1~1_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000000000000110000000011001111000000001100111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_vAluSrc1~2_combout\,
	datac => \ALT_INV_R.curPC\(25),
	datad => \ALT_INV_vAluSrc1~1_combout\,
	dataf => \ALT_INV_Mux65~13_combout\,
	combout => \Mux229~0_combout\);

-- Location: FF_X74_Y3_N40
\R.aluData1[25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux229~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData1\(25));

-- Location: MLABCELL_X78_Y5_N21
\Add1~109\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~109_sumout\ = SUM(( \R.aluData2\(27) ) + ( \R.aluData1\(27) ) + ( \Add1~106\ ))
-- \Add1~110\ = CARRY(( \R.aluData2\(27) ) + ( \R.aluData1\(27) ) + ( \Add1~106\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(27),
	datac => \ALT_INV_R.aluData1\(27),
	cin => \Add1~106\,
	sumout => \Add1~109_sumout\,
	cout => \Add1~110\);

-- Location: MLABCELL_X78_Y5_N24
\Add1~113\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~113_sumout\ = SUM(( \R.aluData2\(28) ) + ( \R.aluData1\(28) ) + ( \Add1~110\ ))
-- \Add1~114\ = CARRY(( \R.aluData2\(28) ) + ( \R.aluData1\(28) ) + ( \Add1~110\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluData1\(28),
	datad => \ALT_INV_R.aluData2\(28),
	cin => \Add1~110\,
	sumout => \Add1~113_sumout\,
	cout => \Add1~114\);

-- Location: MLABCELL_X82_Y4_N15
\Selector3~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector3~3_combout\ = ( \Add1~117_sumout\ & ( \Add2~117_sumout\ & ( ((\Selector3~2_combout\) # (\R.aluOp.ALUOpSub~q\)) # (\R.aluOp.ALUOpAdd~q\) ) ) ) # ( !\Add1~117_sumout\ & ( \Add2~117_sumout\ & ( (\Selector3~2_combout\) # (\R.aluOp.ALUOpSub~q\) ) ) ) 
-- # ( \Add1~117_sumout\ & ( !\Add2~117_sumout\ & ( (\Selector3~2_combout\) # (\R.aluOp.ALUOpAdd~q\) ) ) ) # ( !\Add1~117_sumout\ & ( !\Add2~117_sumout\ & ( \Selector3~2_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111010111110101111100111111001111110111111101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_Selector3~2_combout\,
	datae => \ALT_INV_Add1~117_sumout\,
	dataf => \ALT_INV_Add2~117_sumout\,
	combout => \Selector3~3_combout\);

-- Location: FF_X82_Y4_N17
\R.aluRes[29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector3~3_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(29));

-- Location: IOIBUF_X20_Y0_N18
\avm_d_readdata[5]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(5),
	o => \avm_d_readdata[5]~input_o\);

-- Location: LABCELL_X79_Y2_N39
\Comb:vRegWriteData[29]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[29]~1_combout\ = ( \avm_d_readdata[23]~input_o\ & ( \avm_d_readdata[5]~input_o\ & ( (!\R.curInst\(14) & ((!\R.curInst\(12) & ((\R.curInst\(13)) # (\avm_d_readdata[31]~input_o\))) # (\R.curInst\(12) & ((!\R.curInst\(13)))))) ) ) ) # ( 
-- !\avm_d_readdata[23]~input_o\ & ( \avm_d_readdata[5]~input_o\ & ( (!\R.curInst\(12) & (!\R.curInst\(14) & ((\R.curInst\(13)) # (\avm_d_readdata[31]~input_o\)))) ) ) ) # ( \avm_d_readdata[23]~input_o\ & ( !\avm_d_readdata[5]~input_o\ & ( (!\R.curInst\(14) 
-- & (!\R.curInst\(13) & ((\avm_d_readdata[31]~input_o\) # (\R.curInst\(12))))) ) ) ) # ( !\avm_d_readdata[23]~input_o\ & ( !\avm_d_readdata[5]~input_o\ & ( (!\R.curInst\(12) & (!\R.curInst\(14) & (\avm_d_readdata[31]~input_o\ & !\R.curInst\(13)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000100000000000010011000000000000001000100010000100110010001000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(12),
	datab => \ALT_INV_R.curInst\(14),
	datac => \ALT_INV_avm_d_readdata[31]~input_o\,
	datad => \ALT_INV_R.curInst\(13),
	datae => \ALT_INV_avm_d_readdata[23]~input_o\,
	dataf => \ALT_INV_avm_d_readdata[5]~input_o\,
	combout => \Comb:vRegWriteData[29]~1_combout\);

-- Location: MLABCELL_X82_Y5_N30
\Comb:vRegWriteData[29]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[29]~2_combout\ = ( \Add1~117_sumout\ & ( \Comb:vRegWriteData[29]~1_combout\ & ( (!\R.memToReg~q\ & (!\Selector3~2_combout\ & !\R.aluOp.ALUOpAdd~q\)) ) ) ) # ( !\Add1~117_sumout\ & ( \Comb:vRegWriteData[29]~1_combout\ & ( 
-- (!\R.memToReg~q\ & !\Selector3~2_combout\) ) ) ) # ( \Add1~117_sumout\ & ( !\Comb:vRegWriteData[29]~1_combout\ & ( ((!\Selector3~2_combout\ & !\R.aluOp.ALUOpAdd~q\)) # (\R.memToReg~q\) ) ) ) # ( !\Add1~117_sumout\ & ( !\Comb:vRegWriteData[29]~1_combout\ & 
-- ( (!\Selector3~2_combout\) # (\R.memToReg~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111001111110011111100110011001111000000110000001100000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.memToReg~q\,
	datac => \ALT_INV_Selector3~2_combout\,
	datad => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datae => \ALT_INV_Add1~117_sumout\,
	dataf => \ALT_INV_Comb:vRegWriteData[29]~1_combout\,
	combout => \Comb:vRegWriteData[29]~2_combout\);

-- Location: MLABCELL_X82_Y5_N48
\Comb:vRegWriteData[29]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[29]~0_combout\ = ( \R.aluOp.ALUOpSub~q\ & ( \Comb:vRegWriteData[29]~2_combout\ & ( (!\R.memToReg~q\ & ((!\R.aluCalc~q\ & (\R.aluRes\(29))) # (\R.aluCalc~q\ & ((\Add2~117_sumout\))))) ) ) ) # ( !\R.aluOp.ALUOpSub~q\ & ( 
-- \Comb:vRegWriteData[29]~2_combout\ & ( (\R.aluRes\(29) & (!\R.memToReg~q\ & !\R.aluCalc~q\)) ) ) ) # ( \R.aluOp.ALUOpSub~q\ & ( !\Comb:vRegWriteData[29]~2_combout\ & ( ((\R.aluCalc~q\) # (\R.memToReg~q\)) # (\R.aluRes\(29)) ) ) ) # ( !\R.aluOp.ALUOpSub~q\ 
-- & ( !\Comb:vRegWriteData[29]~2_combout\ & ( ((\R.aluCalc~q\) # (\R.memToReg~q\)) # (\R.aluRes\(29)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0111111101111111011111110111111101000000010000000100000001001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluRes\(29),
	datab => \ALT_INV_R.memToReg~q\,
	datac => \ALT_INV_R.aluCalc~q\,
	datad => \ALT_INV_Add2~117_sumout\,
	datae => \ALT_INV_R.aluOp.ALUOpSub~q\,
	dataf => \ALT_INV_Comb:vRegWriteData[29]~2_combout\,
	combout => \Comb:vRegWriteData[29]~0_combout\);

-- Location: FF_X81_Y5_N53
\R.regWriteData[29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Add0~109_sumout\,
	asdata => \Comb:vRegWriteData[29]~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(29));

-- Location: FF_X67_Y1_N38
\RegFile[31][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(29),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][29]~q\);

-- Location: LABCELL_X68_Y1_N0
\RegFile[30][29]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[30][29]~feeder_combout\ = ( \R.regWriteData\(29) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(29),
	combout => \RegFile[30][29]~feeder_combout\);

-- Location: FF_X68_Y1_N2
\RegFile[30][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[30][29]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][29]~q\);

-- Location: FF_X68_Y1_N44
\RegFile[29][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(29),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][29]~q\);

-- Location: FF_X67_Y1_N26
\RegFile[27][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(29),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][29]~q\);

-- Location: FF_X67_Y1_N8
\RegFile[25][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(29),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][29]~q\);

-- Location: FF_X60_Y2_N28
\RegFile[26][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(29),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][29]~q\);

-- Location: MLABCELL_X59_Y2_N48
\RegFile[24][29]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[24][29]~feeder_combout\ = ( \R.regWriteData\(29) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(29),
	combout => \RegFile[24][29]~feeder_combout\);

-- Location: FF_X59_Y2_N49
\RegFile[24][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[24][29]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][29]~q\);

-- Location: LABCELL_X67_Y1_N6
\Mux93~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux93~22_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[24][29]~q\))) # (\R.curInst\(20) & (\RegFile[25][29]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[26][29]~q\))) # (\R.curInst\(20) & (\RegFile[27][29]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[27][29]~q\,
	datab => \ALT_INV_RegFile[25][29]~q\,
	datac => \ALT_INV_RegFile[26][29]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][29]~q\,
	combout => \Mux93~22_combout\);

-- Location: LABCELL_X73_Y2_N48
\RegFile[28][29]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[28][29]~feeder_combout\ = ( \R.regWriteData\(29) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(29),
	combout => \RegFile[28][29]~feeder_combout\);

-- Location: FF_X73_Y2_N49
\RegFile[28][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[28][29]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][29]~q\);

-- Location: LABCELL_X68_Y1_N42
\Mux93~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux93~9_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux93~22_combout\)))) # (\R.curInst\(22) & ((!\Mux93~22_combout\ & (\RegFile[28][29]~q\)) # (\Mux93~22_combout\ & ((\RegFile[29][29]~q\)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) 
-- & ((((\Mux93~22_combout\))))) # (\R.curInst\(22) & (((!\Mux93~22_combout\ & ((\RegFile[30][29]~q\))) # (\Mux93~22_combout\ & (\RegFile[31][29]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111001100111111111101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][29]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[30][29]~q\,
	datad => \ALT_INV_RegFile[29][29]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux93~22_combout\,
	datag => \ALT_INV_RegFile[28][29]~q\,
	combout => \Mux93~9_combout\);

-- Location: FF_X65_Y2_N26
\RegFile[23][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(29),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][29]~q\);

-- Location: MLABCELL_X59_Y2_N36
\RegFile[22][29]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[22][29]~feeder_combout\ = ( \R.regWriteData\(29) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(29),
	combout => \RegFile[22][29]~feeder_combout\);

-- Location: FF_X59_Y2_N37
\RegFile[22][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[22][29]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][29]~q\);

-- Location: FF_X71_Y2_N26
\RegFile[21][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(29),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][29]~q\);

-- Location: FF_X65_Y2_N14
\RegFile[19][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(29),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][29]~q\);

-- Location: FF_X65_Y2_N8
\RegFile[17][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(29),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][29]~q\);

-- Location: MLABCELL_X59_Y3_N12
\RegFile[18][29]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[18][29]~feeder_combout\ = ( \R.regWriteData\(29) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(29),
	combout => \RegFile[18][29]~feeder_combout\);

-- Location: FF_X59_Y3_N13
\RegFile[18][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][29]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][29]~q\);

-- Location: FF_X64_Y1_N4
\RegFile[16][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(29),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][29]~q\);

-- Location: MLABCELL_X65_Y2_N6
\Mux93~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux93~18_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[16][29]~q\))) # (\R.curInst\(20) & (\RegFile[17][29]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[18][29]~q\))) # (\R.curInst\(20) & (\RegFile[19][29]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[19][29]~q\,
	datab => \ALT_INV_RegFile[17][29]~q\,
	datac => \ALT_INV_RegFile[18][29]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][29]~q\,
	combout => \Mux93~18_combout\);

-- Location: MLABCELL_X59_Y3_N48
\RegFile[20][29]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[20][29]~feeder_combout\ = ( \R.regWriteData\(29) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(29),
	combout => \RegFile[20][29]~feeder_combout\);

-- Location: FF_X59_Y3_N49
\RegFile[20][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[20][29]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][29]~q\);

-- Location: LABCELL_X71_Y2_N24
\Mux93~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux93~5_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux93~18_combout\))))) # (\R.curInst\(22) & (((!\Mux93~18_combout\ & (\RegFile[20][29]~q\)) # (\Mux93~18_combout\ & ((\RegFile[21][29]~q\)))))) ) ) # ( \R.curInst\(21) & ( 
-- (!\R.curInst\(22) & ((((\Mux93~18_combout\))))) # (\R.curInst\(22) & (((!\Mux93~18_combout\ & ((\RegFile[22][29]~q\))) # (\Mux93~18_combout\ & (\RegFile[23][29]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110101010111111111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[23][29]~q\,
	datac => \ALT_INV_RegFile[22][29]~q\,
	datad => \ALT_INV_RegFile[21][29]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux93~18_combout\,
	datag => \ALT_INV_RegFile[20][29]~q\,
	combout => \Mux93~5_combout\);

-- Location: FF_X67_Y3_N43
\RegFile[3][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(29),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][29]~q\);

-- Location: FF_X68_Y1_N56
\RegFile[2][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(29),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][29]~q\);

-- Location: FF_X67_Y3_N2
\RegFile[7][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(29),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][29]~q\);

-- Location: LABCELL_X60_Y3_N57
\RegFile[4][29]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[4][29]~feeder_combout\ = ( \R.regWriteData\(29) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(29),
	combout => \RegFile[4][29]~feeder_combout\);

-- Location: FF_X60_Y3_N58
\RegFile[4][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[4][29]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][29]~q\);

-- Location: FF_X67_Y3_N11
\RegFile[6][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(29),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][29]~q\);

-- Location: FF_X62_Y3_N28
\RegFile[5][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(29),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][29]~q\);

-- Location: LABCELL_X62_Y3_N27
\Mux93~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux93~0_combout\ = ( \RegFile[5][29]~q\ & ( \R.curInst\(20) & ( (!\R.curInst\(21)) # (\RegFile[7][29]~q\) ) ) ) # ( !\RegFile[5][29]~q\ & ( \R.curInst\(20) & ( (\R.curInst\(21) & \RegFile[7][29]~q\) ) ) ) # ( \RegFile[5][29]~q\ & ( !\R.curInst\(20) & ( 
-- (!\R.curInst\(21) & (\RegFile[4][29]~q\)) # (\R.curInst\(21) & ((\RegFile[6][29]~q\))) ) ) ) # ( !\RegFile[5][29]~q\ & ( !\R.curInst\(20) & ( (!\R.curInst\(21) & (\RegFile[4][29]~q\)) # (\R.curInst\(21) & ((\RegFile[6][29]~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101001011111000010100101111100010001000100011011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(21),
	datab => \ALT_INV_RegFile[7][29]~q\,
	datac => \ALT_INV_RegFile[4][29]~q\,
	datad => \ALT_INV_RegFile[6][29]~q\,
	datae => \ALT_INV_RegFile[5][29]~q\,
	dataf => \ALT_INV_R.curInst\(20),
	combout => \Mux93~0_combout\);

-- Location: FF_X61_Y5_N28
\RegFile[1][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(29),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][29]~q\);

-- Location: LABCELL_X68_Y1_N54
\Mux93~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux93~26_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (\R.curInst\(20) & (\RegFile[1][29]~q\))) # (\R.curInst\(22) & (((\Mux93~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (((\RegFile[2][29]~q\)))) # 
-- (\R.curInst\(20) & (\RegFile[3][29]~q\)))) # (\R.curInst\(22) & ((((\Mux93~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000000000111010000000000000011111111110001110111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][29]~q\,
	datab => \ALT_INV_R.curInst\(20),
	datac => \ALT_INV_RegFile[2][29]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux93~0_combout\,
	datag => \ALT_INV_RegFile[1][29]~q\,
	combout => \Mux93~26_combout\);

-- Location: LABCELL_X71_Y2_N36
\RegFile[13][29]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[13][29]~feeder_combout\ = ( \R.regWriteData\(29) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(29),
	combout => \RegFile[13][29]~feeder_combout\);

-- Location: FF_X71_Y2_N37
\RegFile[13][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[13][29]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][29]~q\);

-- Location: LABCELL_X62_Y2_N18
\RegFile[14][29]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[14][29]~feeder_combout\ = ( \R.regWriteData\(29) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(29),
	combout => \RegFile[14][29]~feeder_combout\);

-- Location: FF_X62_Y2_N19
\RegFile[14][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[14][29]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][29]~q\);

-- Location: FF_X70_Y1_N56
\RegFile[15][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(29),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][29]~q\);

-- Location: FF_X70_Y1_N20
\RegFile[11][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(29),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][29]~q\);

-- Location: LABCELL_X64_Y3_N51
\RegFile[10][29]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[10][29]~feeder_combout\ = \R.regWriteData\(29)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101010101010101010101010101010101010101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.regWriteData\(29),
	combout => \RegFile[10][29]~feeder_combout\);

-- Location: FF_X64_Y3_N52
\RegFile[10][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[10][29]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][29]~q\);

-- Location: FF_X72_Y2_N25
\RegFile[9][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(29),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][29]~q\);

-- Location: FF_X66_Y5_N17
\RegFile[8][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(29),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][29]~q\);

-- Location: LABCELL_X71_Y2_N48
\Mux93~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux93~14_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & (\RegFile[8][29]~q\)) # (\R.curInst\(20) & ((\RegFile[9][29]~q\)))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & ((\RegFile[10][29]~q\))) # (\R.curInst\(20) & (\RegFile[11][29]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001010101111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[11][29]~q\,
	datac => \ALT_INV_RegFile[10][29]~q\,
	datad => \ALT_INV_RegFile[9][29]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][29]~q\,
	combout => \Mux93~14_combout\);

-- Location: FF_X74_Y1_N34
\RegFile[12][29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(29),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][29]~q\);

-- Location: LABCELL_X70_Y1_N15
\Mux93~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux93~1_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux93~14_combout\))))) # (\R.curInst\(22) & (((!\Mux93~14_combout\ & ((\RegFile[12][29]~q\))) # (\Mux93~14_combout\ & (\RegFile[13][29]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux93~14_combout\)))) # (\R.curInst\(22) & ((!\Mux93~14_combout\ & (\RegFile[14][29]~q\)) # (\Mux93~14_combout\ & ((\RegFile[15][29]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][29]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[14][29]~q\,
	datad => \ALT_INV_RegFile[15][29]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux93~14_combout\,
	datag => \ALT_INV_RegFile[12][29]~q\,
	combout => \Mux93~1_combout\);

-- Location: LABCELL_X73_Y1_N39
\Mux93~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux93~13_combout\ = ( \Mux93~26_combout\ & ( \Mux93~1_combout\ & ( (!\R.curInst\(24)) # ((!\R.curInst\(23) & ((\Mux93~5_combout\))) # (\R.curInst\(23) & (\Mux93~9_combout\))) ) ) ) # ( !\Mux93~26_combout\ & ( \Mux93~1_combout\ & ( (!\R.curInst\(24) & 
-- (((\R.curInst\(23))))) # (\R.curInst\(24) & ((!\R.curInst\(23) & ((\Mux93~5_combout\))) # (\R.curInst\(23) & (\Mux93~9_combout\)))) ) ) ) # ( \Mux93~26_combout\ & ( !\Mux93~1_combout\ & ( (!\R.curInst\(24) & (((!\R.curInst\(23))))) # (\R.curInst\(24) & 
-- ((!\R.curInst\(23) & ((\Mux93~5_combout\))) # (\R.curInst\(23) & (\Mux93~9_combout\)))) ) ) ) # ( !\Mux93~26_combout\ & ( !\Mux93~1_combout\ & ( (\R.curInst\(24) & ((!\R.curInst\(23) & ((\Mux93~5_combout\))) # (\R.curInst\(23) & (\Mux93~9_combout\)))) ) ) 
-- )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000101010001101000011111000100001011010110111010101111111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(24),
	datab => \ALT_INV_Mux93~9_combout\,
	datac => \ALT_INV_R.curInst\(23),
	datad => \ALT_INV_Mux93~5_combout\,
	datae => \ALT_INV_Mux93~26_combout\,
	dataf => \ALT_INV_Mux93~1_combout\,
	combout => \Mux93~13_combout\);

-- Location: LABCELL_X75_Y3_N36
\NxR.aluData2[29]~31\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[29]~31_combout\ = ( \Mux125~0_combout\ & ( \Mux93~13_combout\ & ( (!\vAluSrc2~1_combout\) # (\Equal4~1_combout\) ) ) ) # ( !\Mux125~0_combout\ & ( \Mux93~13_combout\ & ( !\vAluSrc2~1_combout\ ) ) ) # ( \Mux125~0_combout\ & ( 
-- !\Mux93~13_combout\ & ( (\Equal4~1_combout\ & \vAluSrc2~1_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000001010000010111110000111100001111010111110101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Equal4~1_combout\,
	datac => \ALT_INV_vAluSrc2~1_combout\,
	datae => \ALT_INV_Mux125~0_combout\,
	dataf => \ALT_INV_Mux93~13_combout\,
	combout => \NxR.aluData2[29]~31_combout\);

-- Location: FF_X75_Y3_N37
\R.aluData2[29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR.aluData2[29]~31_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData2\(29));

-- Location: MLABCELL_X82_Y4_N24
\Selector3~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector3~1_combout\ = ( \R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( \R.aluOp.ALUOpOr~q\ & ( (!\R.aluData1\(29) & (!\Selector17~0_OTERM391\ & !\R.aluData2\(29))) ) ) ) # ( !\R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( \R.aluOp.ALUOpOr~q\ & ( (!\R.aluData1\(29) & 
-- (!\Selector17~0_OTERM391\ & !\R.aluData2\(29))) ) ) ) # ( \R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( !\R.aluOp.ALUOpOr~q\ & ( (!\Selector17~0_OTERM391\ & ((!\R.aluOp.ALUOpXor~DUPLICATE_q\ & ((!\R.aluData1\(29)) # (!\R.aluData2\(29)))) # 
-- (\R.aluOp.ALUOpXor~DUPLICATE_q\ & (!\R.aluData1\(29) & !\R.aluData2\(29))))) ) ) ) # ( !\R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( !\R.aluOp.ALUOpOr~q\ & ( (!\Selector17~0_OTERM391\ & ((!\R.aluOp.ALUOpXor~DUPLICATE_q\) # (!\R.aluData1\(29) $ (\R.aluData2\(29))))) 
-- ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1110000010110000111000001000000011000000000000001100000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpXor~DUPLICATE_q\,
	datab => \ALT_INV_R.aluData1\(29),
	datac => \ALT_INV_Selector17~0_OTERM391\,
	datad => \ALT_INV_R.aluData2\(29),
	datae => \ALT_INV_R.aluOp.ALUOpAnd~DUPLICATE_q\,
	dataf => \ALT_INV_R.aluOp.ALUOpOr~q\,
	combout => \Selector3~1_combout\);

-- Location: LABCELL_X80_Y7_N6
\ShiftLeft0~19\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~19_combout\ = ( \ShiftLeft0~1_OTERM255\ & ( \ShiftLeft0~18_OTERM289\ & ( (!\R.aluData2\(3) & ((!\R.aluData2\(2)) # ((\ShiftLeft0~12_OTERM791\)))) # (\R.aluData2\(3) & (((\ShiftLeft0~7_OTERM205\)) # (\R.aluData2\(2)))) ) ) ) # ( 
-- !\ShiftLeft0~1_OTERM255\ & ( \ShiftLeft0~18_OTERM289\ & ( (!\R.aluData2\(3) & ((!\R.aluData2\(2)) # ((\ShiftLeft0~12_OTERM791\)))) # (\R.aluData2\(3) & (!\R.aluData2\(2) & ((\ShiftLeft0~7_OTERM205\)))) ) ) ) # ( \ShiftLeft0~1_OTERM255\ & ( 
-- !\ShiftLeft0~18_OTERM289\ & ( (!\R.aluData2\(3) & (\R.aluData2\(2) & (\ShiftLeft0~12_OTERM791\))) # (\R.aluData2\(3) & (((\ShiftLeft0~7_OTERM205\)) # (\R.aluData2\(2)))) ) ) ) # ( !\ShiftLeft0~1_OTERM255\ & ( !\ShiftLeft0~18_OTERM289\ & ( 
-- (!\R.aluData2\(3) & (\R.aluData2\(2) & (\ShiftLeft0~12_OTERM791\))) # (\R.aluData2\(3) & (!\R.aluData2\(2) & ((\ShiftLeft0~7_OTERM205\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001001000110000100110101011110001010110011101001101111011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(3),
	datab => \ALT_INV_R.aluData2\(2),
	datac => \ALT_INV_ShiftLeft0~12_OTERM791\,
	datad => \ALT_INV_ShiftLeft0~7_OTERM205\,
	datae => \ALT_INV_ShiftLeft0~1_OTERM255\,
	dataf => \ALT_INV_ShiftLeft0~18_OTERM289\,
	combout => \ShiftLeft0~19_combout\);

-- Location: LABCELL_X73_Y5_N18
\ShiftLeft0~51\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~51_combout\ = ( \Mux227~0_combout\ & ( \NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (\Mux226~0_combout\)) # (\NxR.aluData2[1]~17_combout\ & ((\Mux228~0_combout\))) ) ) ) # ( !\Mux227~0_combout\ & ( 
-- \NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (\Mux226~0_combout\)) # (\NxR.aluData2[1]~17_combout\ & ((\Mux228~0_combout\))) ) ) ) # ( \Mux227~0_combout\ & ( !\NxR.aluData2[0]~16_combout\ & ( (\NxR.aluData2[1]~17_combout\) # 
-- (\Mux225~0_combout\) ) ) ) # ( !\Mux227~0_combout\ & ( !\NxR.aluData2[0]~16_combout\ & ( (\Mux225~0_combout\ & !\NxR.aluData2[1]~17_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100010001000100011101110111011100001100001111110000110000111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux225~0_combout\,
	datab => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datac => \ALT_INV_Mux226~0_combout\,
	datad => \ALT_INV_Mux228~0_combout\,
	datae => \ALT_INV_Mux227~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[0]~16_combout\,
	combout => \ShiftLeft0~51_combout\);

-- Location: FF_X73_Y5_N19
\ShiftLeft0~51_NEW_REG762\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~51_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~51_OTERM763\);

-- Location: LABCELL_X83_Y4_N48
\ShiftLeft0~52\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~52_combout\ = ( \R.aluData2\(3) & ( \ShiftLeft0~26_OTERM739\ & ( (\ShiftLeft0~34_OTERM299\) # (\R.aluData2\(2)) ) ) ) # ( !\R.aluData2\(3) & ( \ShiftLeft0~26_OTERM739\ & ( (!\R.aluData2\(2) & (\ShiftLeft0~51_OTERM763\)) # (\R.aluData2\(2) & 
-- ((\ShiftLeft0~42_OTERM41\))) ) ) ) # ( \R.aluData2\(3) & ( !\ShiftLeft0~26_OTERM739\ & ( (!\R.aluData2\(2) & \ShiftLeft0~34_OTERM299\) ) ) ) # ( !\R.aluData2\(3) & ( !\ShiftLeft0~26_OTERM739\ & ( (!\R.aluData2\(2) & (\ShiftLeft0~51_OTERM763\)) # 
-- (\R.aluData2\(2) & ((\ShiftLeft0~42_OTERM41\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101001011111001000100010001000001010010111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(2),
	datab => \ALT_INV_ShiftLeft0~34_OTERM299\,
	datac => \ALT_INV_ShiftLeft0~51_OTERM763\,
	datad => \ALT_INV_ShiftLeft0~42_OTERM41\,
	datae => \ALT_INV_R.aluData2\(3),
	dataf => \ALT_INV_ShiftLeft0~26_OTERM739\,
	combout => \ShiftLeft0~52_combout\);

-- Location: MLABCELL_X82_Y5_N45
\Selector3~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector3~0_combout\ = ( \ShiftRight0~7_OTERM233DUPLICATE_q\ & ( \R.aluData1\(31) & ( \R.aluOp.ALUOpSRA~q\ ) ) ) # ( !\ShiftRight0~7_OTERM233DUPLICATE_q\ & ( \R.aluData1\(31) & ( (!\R.aluOp.ALUOpSRL~q\ & (((\R.aluOp.ALUOpSRA~q\ & 
-- \ShiftRight1~13_OTERM15\)))) # (\R.aluOp.ALUOpSRL~q\ & (((\R.aluOp.ALUOpSRA~q\ & \ShiftRight1~13_OTERM15\)) # (\ShiftRight0~0_OTERM17\))) ) ) ) # ( !\ShiftRight0~7_OTERM233DUPLICATE_q\ & ( !\R.aluData1\(31) & ( (!\R.aluOp.ALUOpSRL~q\ & 
-- (((\R.aluOp.ALUOpSRA~q\ & \ShiftRight1~13_OTERM15\)))) # (\R.aluOp.ALUOpSRL~q\ & (((\R.aluOp.ALUOpSRA~q\ & \ShiftRight1~13_OTERM15\)) # (\ShiftRight0~0_OTERM17\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100011111000000000000000000010001000111110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpSRL~q\,
	datab => \ALT_INV_ShiftRight0~0_OTERM17\,
	datac => \ALT_INV_R.aluOp.ALUOpSRA~q\,
	datad => \ALT_INV_ShiftRight1~13_OTERM15\,
	datae => \ALT_INV_ShiftRight0~7_OTERM233DUPLICATE_q\,
	dataf => \ALT_INV_R.aluData1\(31),
	combout => \Selector3~0_combout\);

-- Location: MLABCELL_X82_Y4_N30
\Selector3~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector3~2_combout\ = ( \ShiftLeft0~52_combout\ & ( \Selector3~0_combout\ & ( (!\Selector3~1_combout\) # ((!\R.aluData2\(4)) # ((\ShiftLeft0~19_combout\ & \R.aluOp.ALUOpSLL~q\))) ) ) ) # ( !\ShiftLeft0~52_combout\ & ( \Selector3~0_combout\ & ( 
-- (!\Selector3~1_combout\) # ((!\R.aluData2\(4)) # ((\ShiftLeft0~19_combout\ & \R.aluOp.ALUOpSLL~q\))) ) ) ) # ( \ShiftLeft0~52_combout\ & ( !\Selector3~0_combout\ & ( (!\Selector3~1_combout\) # ((\R.aluOp.ALUOpSLL~q\ & ((!\R.aluData2\(4)) # 
-- (\ShiftLeft0~19_combout\)))) ) ) ) # ( !\ShiftLeft0~52_combout\ & ( !\Selector3~0_combout\ & ( (!\Selector3~1_combout\) # ((\ShiftLeft0~19_combout\ & (\R.aluData2\(4) & \R.aluOp.ALUOpSLL~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010101010101011101010101111101111111010111110111111101011111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector3~1_combout\,
	datab => \ALT_INV_ShiftLeft0~19_combout\,
	datac => \ALT_INV_R.aluData2\(4),
	datad => \ALT_INV_R.aluOp.ALUOpSLL~q\,
	datae => \ALT_INV_ShiftLeft0~52_combout\,
	dataf => \ALT_INV_Selector3~0_combout\,
	combout => \Selector3~2_combout\);

-- Location: LABCELL_X79_Y4_N42
\Comb:vJumpAdr[29]~0_RESYN1034\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[29]~0_RESYN1034_BDD1035\ = ( \Add2~117_sumout\ & ( ((\R.aluOp.ALUOpAdd~q\ & \Add1~117_sumout\)) # (\R.aluOp.ALUOpSub~q\) ) ) # ( !\Add2~117_sumout\ & ( (\R.aluOp.ALUOpAdd~q\ & \Add1~117_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010101000000000101010100001111010111110000111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datac => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datad => \ALT_INV_Add1~117_sumout\,
	dataf => \ALT_INV_Add2~117_sumout\,
	combout => \Comb:vJumpAdr[29]~0_RESYN1034_BDD1035\);

-- Location: LABCELL_X74_Y4_N42
\Mux126~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux126~0_combout\ = ( \R.curInst\(28) & ( ((\vAluSrc1~0_combout\ & ((\R.curInst\(2)) # (\Mux124~0_combout\)))) # (\Mux123~1_combout\) ) ) # ( !\R.curInst\(28) & ( ((\Mux124~0_combout\ & \vAluSrc1~0_combout\)) # (\Mux123~1_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010111111111000001011111111100000111111111110000011111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux124~0_combout\,
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_vAluSrc1~0_combout\,
	datad => \ALT_INV_Mux123~1_combout\,
	dataf => \ALT_INV_R.curInst\(28),
	combout => \Mux126~0_combout\);

-- Location: LABCELL_X75_Y4_N9
\Mux133~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux133~0_combout\ = ( \R.curInst\(21) & ( ((\vAluSrc1~0_combout\ & ((\Mux124~0_combout\) # (\R.curInst\(2))))) # (\Mux123~1_combout\) ) ) # ( !\R.curInst\(21) & ( ((\vAluSrc1~0_combout\ & \Mux124~0_combout\)) # (\Mux123~1_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111101011111000011110101111100011111010111110001111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluSrc1~0_combout\,
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_Mux123~1_combout\,
	datad => \ALT_INV_Mux124~0_combout\,
	dataf => \ALT_INV_R.curInst\(21),
	combout => \Mux133~0_combout\);

-- Location: FF_X78_Y2_N35
\R.curPC[21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[21]~0_combout\,
	asdata => \Add0~77_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(21));

-- Location: LABCELL_X77_Y4_N27
\Add3~77\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~77_sumout\ = SUM(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux135~0_combout\)) ) + ( \R.curPC\(19) ) + ( \Add3~74\ ))
-- \Add3~78\ = CARRY(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux135~0_combout\)) ) + ( \R.curPC\(19) ) + ( \Add3~74\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000010001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datac => \ALT_INV_R.curPC\(19),
	datad => \ALT_INV_Mux135~0_combout\,
	cin => \Add3~74\,
	sumout => \Add3~77_sumout\,
	cout => \Add3~78\);

-- Location: LABCELL_X77_Y4_N30
\Add3~81\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~81_sumout\ = SUM(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux134~0_combout\)) ) + ( \R.curPC\(20) ) + ( \Add3~78\ ))
-- \Add3~82\ = CARRY(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux134~0_combout\)) ) + ( \R.curPC\(20) ) + ( \Add3~78\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000000000010001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datad => \ALT_INV_Mux134~0_combout\,
	dataf => \ALT_INV_R.curPC\(20),
	cin => \Add3~78\,
	sumout => \Add3~81_sumout\,
	cout => \Add3~82\);

-- Location: LABCELL_X77_Y4_N33
\Add3~85\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~85_sumout\ = SUM(( \R.curPC\(21) ) + ( (\R.curInst\(0) & (\R.curInst\(1) & \Mux133~0_combout\)) ) + ( \Add3~82\ ))
-- \Add3~86\ = CARRY(( \R.curPC\(21) ) + ( (\R.curInst\(0) & (\R.curInst\(1) & \Mux133~0_combout\)) ) + ( \Add3~82\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111101111111000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datac => \ALT_INV_Mux133~0_combout\,
	datad => \ALT_INV_R.curPC\(21),
	cin => \Add3~82\,
	sumout => \Add3~85_sumout\,
	cout => \Add3~86\);

-- Location: LABCELL_X77_Y4_N36
\Add3~89\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~89_sumout\ = SUM(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux132~0_combout\)) ) + ( \R.curPC\(22) ) + ( \Add3~86\ ))
-- \Add3~90\ = CARRY(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux132~0_combout\)) ) + ( \R.curPC\(22) ) + ( \Add3~86\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000000000010001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datad => \ALT_INV_Mux132~0_combout\,
	dataf => \ALT_INV_R.curPC\(22),
	cin => \Add3~86\,
	sumout => \Add3~89_sumout\,
	cout => \Add3~90\);

-- Location: LABCELL_X77_Y4_N39
\Add3~93\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~93_sumout\ = SUM(( \R.curPC\(23) ) + ( (\R.curInst\(0) & (\R.curInst\(1) & \Mux131~0_combout\)) ) + ( \Add3~90\ ))
-- \Add3~94\ = CARRY(( \R.curPC\(23) ) + ( (\R.curInst\(0) & (\R.curInst\(1) & \Mux131~0_combout\)) ) + ( \Add3~90\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111101111111000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datac => \ALT_INV_Mux131~0_combout\,
	datad => \ALT_INV_R.curPC\(23),
	cin => \Add3~90\,
	sumout => \Add3~93_sumout\,
	cout => \Add3~94\);

-- Location: LABCELL_X77_Y4_N42
\Add3~97\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~97_sumout\ = SUM(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux130~0_combout\)) ) + ( \R.curPC\(24) ) + ( \Add3~94\ ))
-- \Add3~98\ = CARRY(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux130~0_combout\)) ) + ( \R.curPC\(24) ) + ( \Add3~94\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000000000010001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datad => \ALT_INV_Mux130~0_combout\,
	dataf => \ALT_INV_R.curPC\(24),
	cin => \Add3~94\,
	sumout => \Add3~97_sumout\,
	cout => \Add3~98\);

-- Location: LABCELL_X77_Y4_N45
\Add3~101\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~101_sumout\ = SUM(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux129~0_combout\)) ) + ( \R.curPC\(25) ) + ( \Add3~98\ ))
-- \Add3~102\ = CARRY(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux129~0_combout\)) ) + ( \R.curPC\(25) ) + ( \Add3~98\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000010001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datac => \ALT_INV_R.curPC\(25),
	datad => \ALT_INV_Mux129~0_combout\,
	cin => \Add3~98\,
	sumout => \Add3~101_sumout\,
	cout => \Add3~102\);

-- Location: LABCELL_X77_Y4_N48
\Add3~105\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~105_sumout\ = SUM(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux128~0_combout\)) ) + ( \R.curPC\(26) ) + ( \Add3~102\ ))
-- \Add3~106\ = CARRY(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux128~0_combout\)) ) + ( \R.curPC\(26) ) + ( \Add3~102\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000010001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datac => \ALT_INV_R.curPC\(26),
	datad => \ALT_INV_Mux128~0_combout\,
	cin => \Add3~102\,
	sumout => \Add3~105_sumout\,
	cout => \Add3~106\);

-- Location: LABCELL_X77_Y4_N51
\Add3~109\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~109_sumout\ = SUM(( \R.curPC\(27) ) + ( (\R.curInst\(0) & (\R.curInst\(1) & \Mux127~0_combout\)) ) + ( \Add3~106\ ))
-- \Add3~110\ = CARRY(( \R.curPC\(27) ) + ( (\R.curInst\(0) & (\R.curInst\(1) & \Mux127~0_combout\)) ) + ( \Add3~106\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111101111111000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datac => \ALT_INV_Mux127~0_combout\,
	datad => \ALT_INV_R.curPC\(27),
	cin => \Add3~106\,
	sumout => \Add3~109_sumout\,
	cout => \Add3~110\);

-- Location: LABCELL_X77_Y4_N54
\Add3~113\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~113_sumout\ = SUM(( \R.curPC\(28) ) + ( (\R.curInst\(0) & (\R.curInst\(1) & \Mux126~0_combout\)) ) + ( \Add3~110\ ))
-- \Add3~114\ = CARRY(( \R.curPC\(28) ) + ( (\R.curInst\(0) & (\R.curInst\(1) & \Mux126~0_combout\)) ) + ( \Add3~110\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111101111111000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datac => \ALT_INV_Mux126~0_combout\,
	datad => \ALT_INV_R.curPC\(28),
	cin => \Add3~110\,
	sumout => \Add3~113_sumout\,
	cout => \Add3~114\);

-- Location: LABCELL_X77_Y4_N57
\Add3~117\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~117_sumout\ = SUM(( \R.curPC\(29) ) + ( (\R.curInst\(0) & (\R.curInst\(1) & \Mux125~0_combout\)) ) + ( \Add3~114\ ))
-- \Add3~118\ = CARRY(( \R.curPC\(29) ) + ( (\R.curInst\(0) & (\R.curInst\(1) & \Mux125~0_combout\)) ) + ( \Add3~114\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111101111111000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datac => \ALT_INV_Mux125~0_combout\,
	datad => \ALT_INV_R.curPC\(29),
	cin => \Add3~114\,
	sumout => \Add3~117_sumout\,
	cout => \Add3~118\);

-- Location: MLABCELL_X78_Y4_N12
\Comb:vJumpAdr[29]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[29]~0_combout\ = ( \Equal4~2_combout\ & ( \Add3~117_sumout\ & ( (!\R.aluCalc~q\ & (((\R.aluRes\(29))))) # (\R.aluCalc~q\ & (((\Comb:vJumpAdr[29]~0_RESYN1034_BDD1035\)) # (\Selector3~2_combout\))) ) ) ) # ( !\Equal4~2_combout\ & ( 
-- \Add3~117_sumout\ ) ) # ( \Equal4~2_combout\ & ( !\Add3~117_sumout\ & ( (!\R.aluCalc~q\ & (((\R.aluRes\(29))))) # (\R.aluCalc~q\ & (((\Comb:vJumpAdr[29]~0_RESYN1034_BDD1035\)) # (\Selector3~2_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000001101010011111111111111111111110011010100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector3~2_combout\,
	datab => \ALT_INV_R.aluRes\(29),
	datac => \ALT_INV_R.aluCalc~q\,
	datad => \ALT_INV_Comb:vJumpAdr[29]~0_RESYN1034_BDD1035\,
	datae => \ALT_INV_Equal4~2_combout\,
	dataf => \ALT_INV_Add3~117_sumout\,
	combout => \Comb:vJumpAdr[29]~0_combout\);

-- Location: FF_X78_Y4_N13
\R.curPC[29]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[29]~0_combout\,
	asdata => \Add0~109_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(29));

-- Location: LABCELL_X67_Y1_N24
\Mux61~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux61~22_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[24][29]~q\))) # (\R.curInst\(15) & (\RegFile[25][29]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[26][29]~q\))) # (\R.curInst\(15) & (\RegFile[27][29]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[27][29]~q\,
	datab => \ALT_INV_RegFile[25][29]~q\,
	datac => \ALT_INV_RegFile[26][29]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][29]~q\,
	combout => \Mux61~22_combout\);

-- Location: LABCELL_X67_Y1_N36
\Mux61~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux61~9_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux61~22_combout\))))) # (\R.curInst\(17) & (((!\Mux61~22_combout\ & ((\RegFile[28][29]~q\))) # (\Mux61~22_combout\ & (\RegFile[29][29]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux61~22_combout\)))) # (\R.curInst\(17) & ((!\Mux61~22_combout\ & (\RegFile[30][29]~q\)) # (\Mux61~22_combout\ & ((\RegFile[31][29]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[29][29]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[30][29]~q\,
	datad => \ALT_INV_RegFile[31][29]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux61~22_combout\,
	datag => \ALT_INV_RegFile[28][29]~q\,
	combout => \Mux61~9_combout\);

-- Location: MLABCELL_X65_Y2_N12
\Mux61~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux61~18_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[16][29]~q\))) # (\R.curInst\(15) & (\RegFile[17][29]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[18][29]~q\))) # (\R.curInst\(15) & (\RegFile[19][29]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[19][29]~q\,
	datab => \ALT_INV_RegFile[17][29]~q\,
	datac => \ALT_INV_RegFile[18][29]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][29]~q\,
	combout => \Mux61~18_combout\);

-- Location: MLABCELL_X65_Y2_N24
\Mux61~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux61~5_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux61~18_combout\)))) # (\R.curInst\(17) & ((!\Mux61~18_combout\ & ((\RegFile[20][29]~q\))) # (\Mux61~18_combout\ & (\RegFile[21][29]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux61~18_combout\)))) # (\R.curInst\(17) & ((!\Mux61~18_combout\ & ((\RegFile[22][29]~q\))) # (\Mux61~18_combout\ & (\RegFile[23][29]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[23][29]~q\,
	datab => \ALT_INV_RegFile[21][29]~q\,
	datac => \ALT_INV_RegFile[22][29]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux61~18_combout\,
	datag => \ALT_INV_RegFile[20][29]~q\,
	combout => \Mux61~5_combout\);

-- Location: LABCELL_X70_Y1_N18
\Mux61~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux61~14_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[8][29]~q\))) # (\R.curInst\(15) & (\RegFile[9][29]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[10][29]~q\))) # (\R.curInst\(15) & (\RegFile[11][29]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[11][29]~q\,
	datab => \ALT_INV_RegFile[9][29]~q\,
	datac => \ALT_INV_RegFile[10][29]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][29]~q\,
	combout => \Mux61~14_combout\);

-- Location: LABCELL_X70_Y1_N54
\Mux61~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux61~1_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux61~14_combout\)))) # (\R.curInst\(17) & ((!\Mux61~14_combout\ & ((\RegFile[12][29]~q\))) # (\Mux61~14_combout\ & (\RegFile[13][29]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux61~14_combout\)))) # (\R.curInst\(17) & ((!\Mux61~14_combout\ & ((\RegFile[14][29]~q\))) # (\Mux61~14_combout\ & (\RegFile[15][29]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][29]~q\,
	datab => \ALT_INV_RegFile[13][29]~q\,
	datac => \ALT_INV_RegFile[14][29]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux61~14_combout\,
	datag => \ALT_INV_RegFile[12][29]~q\,
	combout => \Mux61~1_combout\);

-- Location: LABCELL_X67_Y3_N0
\Mux61~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux61~0_combout\ = ( \RegFile[7][29]~q\ & ( \R.curInst\(15) & ( (\RegFile[5][29]~q\) # (\R.curInst\(16)) ) ) ) # ( !\RegFile[7][29]~q\ & ( \R.curInst\(15) & ( (!\R.curInst\(16) & \RegFile[5][29]~q\) ) ) ) # ( \RegFile[7][29]~q\ & ( !\R.curInst\(15) & ( 
-- (!\R.curInst\(16) & (\RegFile[4][29]~q\)) # (\R.curInst\(16) & ((\RegFile[6][29]~q\))) ) ) ) # ( !\RegFile[7][29]~q\ & ( !\R.curInst\(15) & ( (!\R.curInst\(16) & (\RegFile[4][29]~q\)) # (\R.curInst\(16) & ((\RegFile[6][29]~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101001011111000010100101111100100010001000100111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(16),
	datab => \ALT_INV_RegFile[5][29]~q\,
	datac => \ALT_INV_RegFile[4][29]~q\,
	datad => \ALT_INV_RegFile[6][29]~q\,
	datae => \ALT_INV_RegFile[7][29]~q\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux61~0_combout\);

-- Location: FF_X61_Y5_N29
\RegFile[1][29]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(29),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][29]~DUPLICATE_q\);

-- Location: LABCELL_X68_Y3_N24
\Mux61~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux61~26_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (\R.curInst\(15) & (\RegFile[1][29]~DUPLICATE_q\))) # (\R.curInst\(17) & ((((\Mux61~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & ((!\R.curInst\(15) & (\RegFile[2][29]~q\)) 
-- # (\R.curInst\(15) & (((\RegFile[3][29]~q\)))))) # (\R.curInst\(17) & ((((\Mux61~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001000000010000010000010101001010111010101110101110101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_R.curInst\(15),
	datac => \ALT_INV_RegFile[2][29]~q\,
	datad => \ALT_INV_RegFile[3][29]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux61~0_combout\,
	datag => \ALT_INV_RegFile[1][29]~DUPLICATE_q\,
	combout => \Mux61~26_combout\);

-- Location: LABCELL_X70_Y1_N42
\Mux61~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux61~13_combout\ = ( \Mux61~1_combout\ & ( \Mux61~26_combout\ & ( (!\R.curInst\(19)) # ((!\R.curInst\(18) & ((\Mux61~5_combout\))) # (\R.curInst\(18) & (\Mux61~9_combout\))) ) ) ) # ( !\Mux61~1_combout\ & ( \Mux61~26_combout\ & ( (!\R.curInst\(19) & 
-- (((!\R.curInst\(18))))) # (\R.curInst\(19) & ((!\R.curInst\(18) & ((\Mux61~5_combout\))) # (\R.curInst\(18) & (\Mux61~9_combout\)))) ) ) ) # ( \Mux61~1_combout\ & ( !\Mux61~26_combout\ & ( (!\R.curInst\(19) & (((\R.curInst\(18))))) # (\R.curInst\(19) & 
-- ((!\R.curInst\(18) & ((\Mux61~5_combout\))) # (\R.curInst\(18) & (\Mux61~9_combout\)))) ) ) ) # ( !\Mux61~1_combout\ & ( !\Mux61~26_combout\ & ( (\R.curInst\(19) & ((!\R.curInst\(18) & ((\Mux61~5_combout\))) # (\R.curInst\(18) & (\Mux61~9_combout\)))) ) ) 
-- )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100010001000001011011101110101111000100011010111110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(19),
	datab => \ALT_INV_Mux61~9_combout\,
	datac => \ALT_INV_Mux61~5_combout\,
	datad => \ALT_INV_R.curInst\(18),
	datae => \ALT_INV_Mux61~1_combout\,
	dataf => \ALT_INV_Mux61~26_combout\,
	combout => \Mux61~13_combout\);

-- Location: LABCELL_X73_Y5_N0
\Mux225~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux225~0_combout\ = ( \Mux61~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC\(29)))) ) ) # ( !\Mux61~13_combout\ & ( (\vAluSrc1~2_combout\ & (\R.curPC\(29) & !\vAluSrc1~1_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000000000001010000000010101111000000001010111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluSrc1~2_combout\,
	datac => \ALT_INV_R.curPC\(29),
	datad => \ALT_INV_vAluSrc1~1_combout\,
	dataf => \ALT_INV_Mux61~13_combout\,
	combout => \Mux225~0_combout\);

-- Location: LABCELL_X73_Y5_N42
\ShiftRight1~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~13_combout\ = ( \Mux224~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((\NxR.aluData2[0]~16_combout\)) # (\Mux225~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (((\Mux223~0_combout\)))) ) ) # ( !\Mux224~0_combout\ & ( 
-- (!\NxR.aluData2[1]~17_combout\ & (\Mux225~0_combout\ & ((!\NxR.aluData2[0]~16_combout\)))) # (\NxR.aluData2[1]~17_combout\ & (((\Mux223~0_combout\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101001100000011010100110000001101010011111100110101001111110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux225~0_combout\,
	datab => \ALT_INV_Mux223~0_combout\,
	datac => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datad => \ALT_INV_NxR.aluData2[0]~16_combout\,
	dataf => \ALT_INV_Mux224~0_combout\,
	combout => \ShiftRight1~13_combout\);

-- Location: FF_X73_Y5_N43
\ShiftRight1~13_NEW_REG14\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~13_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~13_OTERM15\);

-- Location: LABCELL_X77_Y9_N18
\ShiftRight1~41\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~41_combout\ = ( \R.aluData2\(3) & ( \ShiftRight1~11_OTERM35\ & ( (!\R.aluData2\(2) & (\ShiftRight1~13_OTERM15\)) # (\R.aluData2\(2) & ((\R.aluData1\(31)))) ) ) ) # ( !\R.aluData2\(3) & ( \ShiftRight1~11_OTERM35\ & ( (!\R.aluData2\(2)) # 
-- (\ShiftRight1~12_OTERM57\) ) ) ) # ( \R.aluData2\(3) & ( !\ShiftRight1~11_OTERM35\ & ( (!\R.aluData2\(2) & (\ShiftRight1~13_OTERM15\)) # (\R.aluData2\(2) & ((\R.aluData1\(31)))) ) ) ) # ( !\R.aluData2\(3) & ( !\ShiftRight1~11_OTERM35\ & ( 
-- (\ShiftRight1~12_OTERM57\ & \R.aluData2\(2)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010101001100110000111111111111010101010011001100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~12_OTERM57\,
	datab => \ALT_INV_ShiftRight1~13_OTERM15\,
	datac => \ALT_INV_R.aluData1\(31),
	datad => \ALT_INV_R.aluData2\(2),
	datae => \ALT_INV_R.aluData2\(3),
	dataf => \ALT_INV_ShiftRight1~11_OTERM35\,
	combout => \ShiftRight1~41_combout\);

-- Location: MLABCELL_X82_Y7_N18
\Selector27~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector27~5_combout\ = ( \Selector27~1_combout\ ) # ( !\Selector27~1_combout\ & ( (!\Selector27~4_combout\) # ((\Selector31~6_OTERM381\ & \ShiftRight1~41_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111100000101111111110000010111111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector31~6_OTERM381\,
	datac => \ALT_INV_ShiftRight1~41_combout\,
	datad => \ALT_INV_Selector27~4_combout\,
	dataf => \ALT_INV_Selector27~1_combout\,
	combout => \Selector27~5_combout\);

-- Location: FF_X82_Y7_N19
\R.aluRes[5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector27~5_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(5));

-- Location: LABCELL_X80_Y8_N27
\vAluRes~5_RESYN1070\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~5_RESYN1070_BDD1071\ = ( \Add2~21_sumout\ & ( ((\ShiftRight1~41_combout\ & \Selector31~6_OTERM381\)) # (\R.aluOp.ALUOpSub~q\) ) ) # ( !\Add2~21_sumout\ & ( (\ShiftRight1~41_combout\ & \Selector31~6_OTERM381\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110011000000000011001100001111001111110000111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_ShiftRight1~41_combout\,
	datac => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datad => \ALT_INV_Selector31~6_OTERM381\,
	dataf => \ALT_INV_Add2~21_sumout\,
	combout => \vAluRes~5_RESYN1070_BDD1071\);

-- Location: MLABCELL_X82_Y8_N39
\vAluRes~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~5_combout\ = ( \Add1~21_sumout\ & ( \vAluRes~5_RESYN1070_BDD1071\ & ( (\R.aluRes\(5)) # (\R.aluCalc~q\) ) ) ) # ( !\Add1~21_sumout\ & ( \vAluRes~5_RESYN1070_BDD1071\ & ( (\R.aluRes\(5)) # (\R.aluCalc~q\) ) ) ) # ( \Add1~21_sumout\ & ( 
-- !\vAluRes~5_RESYN1070_BDD1071\ & ( (!\R.aluCalc~q\ & (((\R.aluRes\(5))))) # (\R.aluCalc~q\ & (((!\Selector27~4_combout\)) # (\R.aluOp.ALUOpAdd~q\))) ) ) ) # ( !\Add1~21_sumout\ & ( !\vAluRes~5_RESYN1070_BDD1071\ & ( (!\R.aluCalc~q\ & (\R.aluRes\(5))) # 
-- (\R.aluCalc~q\ & ((!\Selector27~4_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101111100001010010111110001101101011111010111110101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluCalc~q\,
	datab => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datac => \ALT_INV_R.aluRes\(5),
	datad => \ALT_INV_Selector27~4_combout\,
	datae => \ALT_INV_Add1~21_sumout\,
	dataf => \ALT_INV_vAluRes~5_RESYN1070_BDD1071\,
	combout => \vAluRes~5_combout\);

-- Location: MLABCELL_X78_Y8_N51
\Comb:vJumpAdr[5]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[5]~0_combout\ = ( \Equal4~2_combout\ & ( \Add3~21_sumout\ & ( \vAluRes~5_combout\ ) ) ) # ( !\Equal4~2_combout\ & ( \Add3~21_sumout\ ) ) # ( \Equal4~2_combout\ & ( !\Add3~21_sumout\ & ( \vAluRes~5_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000111111111111111111110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_vAluRes~5_combout\,
	datae => \ALT_INV_Equal4~2_combout\,
	dataf => \ALT_INV_Add3~21_sumout\,
	combout => \Comb:vJumpAdr[5]~0_combout\);

-- Location: FF_X78_Y8_N52
\R.curPC[5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[5]~0_combout\,
	asdata => \Add0~13_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(5));

-- Location: LABCELL_X81_Y6_N15
\Add0~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~21_sumout\ = SUM(( \R.curPC\(7) ) + ( GND ) + ( \Add0~18\ ))
-- \Add0~22\ = CARRY(( \R.curPC\(7) ) + ( GND ) + ( \Add0~18\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.curPC\(7),
	cin => \Add0~18\,
	sumout => \Add0~21_sumout\,
	cout => \Add0~22\);

-- Location: LABCELL_X83_Y6_N33
\R.regWriteData[7]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.regWriteData[7]~feeder_combout\ = \Add0~21_sumout\

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101010101010101010101010101010101010101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add0~21_sumout\,
	combout => \R.regWriteData[7]~feeder_combout\);

-- Location: MLABCELL_X84_Y4_N42
\vAluRes~7_RESYN1076_RESYN1132\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~7_RESYN1076_RESYN1132_BDD1133\ = ( \R.aluCalc~q\ & ( \R.aluRes\(7) & ( \Selector31~5_OTERM599\ ) ) ) # ( !\R.aluCalc~q\ & ( \R.aluRes\(7) ) ) # ( \R.aluCalc~q\ & ( !\R.aluRes\(7) & ( \Selector31~5_OTERM599\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000001100110011001111111111111111110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Selector31~5_OTERM599\,
	datae => \ALT_INV_R.aluCalc~q\,
	dataf => \ALT_INV_R.aluRes\(7),
	combout => \vAluRes~7_RESYN1076_RESYN1132_BDD1133\);

-- Location: LABCELL_X83_Y5_N36
\vAluRes~7_RESYN1076\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~7_RESYN1076_BDD1077\ = ( \R.aluCalc~q\ & ( \Selector25~2_combout\ ) ) # ( !\R.aluCalc~q\ & ( \Selector25~2_combout\ & ( \vAluRes~7_RESYN1076_RESYN1132_BDD1133\ ) ) ) # ( \R.aluCalc~q\ & ( !\Selector25~2_combout\ & ( (!\Selector25~4_combout\) # 
-- (((\ShiftRight1~45_combout\ & \vAluRes~7_RESYN1076_RESYN1132_BDD1133\)) # (\Selector25~1_combout\)) ) ) ) # ( !\R.aluCalc~q\ & ( !\Selector25~2_combout\ & ( \vAluRes~7_RESYN1076_RESYN1132_BDD1133\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111101010111111111100001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector25~4_combout\,
	datab => \ALT_INV_ShiftRight1~45_combout\,
	datac => \ALT_INV_vAluRes~7_RESYN1076_RESYN1132_BDD1133\,
	datad => \ALT_INV_Selector25~1_combout\,
	datae => \ALT_INV_R.aluCalc~q\,
	dataf => \ALT_INV_Selector25~2_combout\,
	combout => \vAluRes~7_RESYN1076_BDD1077\);

-- Location: LABCELL_X83_Y5_N12
\Comb:vRegWriteData[7]~0_RESYN1118\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[7]~0_RESYN1118_BDD1119\ = ( \Add2~29_sumout\ & ( (!\R.memToReg~q\ & (((\R.aluOp.ALUOpSub~q\)))) # (\R.memToReg~q\ & (\Mux222~0_combout\ & (\avm_d_readdata[31]~input_o\))) ) ) # ( !\Add2~29_sumout\ & ( (\R.memToReg~q\ & 
-- (\Mux222~0_combout\ & \avm_d_readdata[31]~input_o\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000100000001000000010000000100000001101010110000000110101011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.memToReg~q\,
	datab => \ALT_INV_Mux222~0_combout\,
	datac => \ALT_INV_avm_d_readdata[31]~input_o\,
	datad => \ALT_INV_R.aluOp.ALUOpSub~q\,
	dataf => \ALT_INV_Add2~29_sumout\,
	combout => \Comb:vRegWriteData[7]~0_RESYN1118_BDD1119\);

-- Location: LABCELL_X83_Y5_N30
\Comb:vRegWriteData[7]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[7]~0_combout\ = ( \vAluRes~7_RESYN1076_BDD1077\ & ( \Comb:vRegWriteData[7]~0_RESYN1118_BDD1119\ ) ) # ( !\vAluRes~7_RESYN1076_BDD1077\ & ( \Comb:vRegWriteData[7]~0_RESYN1118_BDD1119\ & ( (\R.aluCalc~q\) # (\R.memToReg~q\) ) ) ) # ( 
-- \vAluRes~7_RESYN1076_BDD1077\ & ( !\Comb:vRegWriteData[7]~0_RESYN1118_BDD1119\ & ( !\R.memToReg~q\ ) ) ) # ( !\vAluRes~7_RESYN1076_BDD1077\ & ( !\Comb:vRegWriteData[7]~0_RESYN1118_BDD1119\ & ( (!\R.memToReg~q\ & (\R.aluCalc~q\ & (\R.aluOp.ALUOpAdd~q\ & 
-- \Add1~29_sumout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000010101010101010101001110111011101111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.memToReg~q\,
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_Add1~29_sumout\,
	datae => \ALT_INV_vAluRes~7_RESYN1076_BDD1077\,
	dataf => \ALT_INV_Comb:vRegWriteData[7]~0_RESYN1118_BDD1119\,
	combout => \Comb:vRegWriteData[7]~0_combout\);

-- Location: FF_X83_Y6_N35
\R.regWriteData[7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \R.regWriteData[7]~feeder_combout\,
	asdata => \Comb:vRegWriteData[7]~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(7));

-- Location: LABCELL_X68_Y7_N54
\RegFile[2][7]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[2][7]~feeder_combout\ = ( \R.regWriteData\(7) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(7),
	combout => \RegFile[2][7]~feeder_combout\);

-- Location: FF_X68_Y7_N56
\RegFile[2][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[2][7]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][7]~q\);

-- Location: LABCELL_X62_Y3_N12
\Mux115~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux115~0_combout\ = ( \RegFile[5][7]~q\ & ( \R.curInst\(20) & ( (!\R.curInst\(21)) # (\RegFile[7][7]~q\) ) ) ) # ( !\RegFile[5][7]~q\ & ( \R.curInst\(20) & ( (\RegFile[7][7]~q\ & \R.curInst\(21)) ) ) ) # ( \RegFile[5][7]~q\ & ( !\R.curInst\(20) & ( 
-- (!\R.curInst\(21) & (\RegFile[4][7]~q\)) # (\R.curInst\(21) & ((\RegFile[6][7]~q\))) ) ) ) # ( !\RegFile[5][7]~q\ & ( !\R.curInst\(20) & ( (!\R.curInst\(21) & (\RegFile[4][7]~q\)) # (\R.curInst\(21) & ((\RegFile[6][7]~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010100110011010101010011001100000000000011111111111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[4][7]~q\,
	datab => \ALT_INV_RegFile[6][7]~q\,
	datac => \ALT_INV_RegFile[7][7]~q\,
	datad => \ALT_INV_R.curInst\(21),
	datae => \ALT_INV_RegFile[5][7]~q\,
	dataf => \ALT_INV_R.curInst\(20),
	combout => \Mux115~0_combout\);

-- Location: LABCELL_X68_Y7_N42
\Mux115~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux115~26_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (\R.curInst\(20) & (\RegFile[1][7]~q\))) # (\R.curInst\(22) & ((((\Mux115~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (\RegFile[2][7]~q\)) # 
-- (\R.curInst\(20) & (((\RegFile[3][7]~q\)))))) # (\R.curInst\(22) & ((((\Mux115~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010000000100000010000100110000110111001101110011101101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(20),
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[2][7]~q\,
	datad => \ALT_INV_RegFile[3][7]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux115~0_combout\,
	datag => \ALT_INV_RegFile[1][7]~q\,
	combout => \Mux115~26_combout\);

-- Location: LABCELL_X63_Y5_N24
\Mux115~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux115~18_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[16][7]~q\))) # (\R.curInst\(20) & (\RegFile[17][7]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[18][7]~q\))) # (\R.curInst\(20) & (\RegFile[19][7]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[17][7]~q\,
	datab => \ALT_INV_RegFile[19][7]~q\,
	datac => \ALT_INV_RegFile[18][7]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][7]~q\,
	combout => \Mux115~18_combout\);

-- Location: LABCELL_X68_Y7_N48
\Mux115~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux115~5_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux115~18_combout\)))) # (\R.curInst\(22) & ((!\Mux115~18_combout\ & ((\RegFile[20][7]~q\))) # (\Mux115~18_combout\ & (\RegFile[21][7]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux115~18_combout\)))) # (\R.curInst\(22) & ((!\Mux115~18_combout\ & ((\RegFile[22][7]~q\))) # (\Mux115~18_combout\ & (\RegFile[23][7]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][7]~q\,
	datab => \ALT_INV_RegFile[23][7]~q\,
	datac => \ALT_INV_RegFile[22][7]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux115~18_combout\,
	datag => \ALT_INV_RegFile[20][7]~q\,
	combout => \Mux115~5_combout\);

-- Location: LABCELL_X61_Y7_N9
\Mux115~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux115~14_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[8][7]~q\))) # (\R.curInst\(20) & (\RegFile[9][7]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & (\RegFile[10][7]~q\)) # (\R.curInst\(20) & ((\RegFile[11][7]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][7]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[10][7]~q\,
	datad => \ALT_INV_RegFile[11][7]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][7]~q\,
	combout => \Mux115~14_combout\);

-- Location: LABCELL_X61_Y7_N24
\Mux115~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux115~1_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux115~14_combout\))))) # (\R.curInst\(22) & (((!\Mux115~14_combout\ & ((\RegFile[12][7]~q\))) # (\Mux115~14_combout\ & (\RegFile[13][7]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux115~14_combout\)))) # (\R.curInst\(22) & ((!\Mux115~14_combout\ & (\RegFile[14][7]~q\)) # (\Mux115~14_combout\ & ((\RegFile[15][7]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][7]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[14][7]~q\,
	datad => \ALT_INV_RegFile[15][7]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux115~14_combout\,
	datag => \ALT_INV_RegFile[12][7]~q\,
	combout => \Mux115~1_combout\);

-- Location: FF_X62_Y6_N7
\RegFile[30][7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[30][7]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][7]~q\);

-- Location: LABCELL_X62_Y4_N30
\Mux115~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux115~22_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[24][7]~q\))) # (\R.curInst\(20) & (\RegFile[25][7]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & (\RegFile[26][7]~q\)) # (\R.curInst\(20) & ((\RegFile[27][7]~q\)))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001110111011101110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[25][7]~q\,
	datac => \ALT_INV_RegFile[26][7]~q\,
	datad => \ALT_INV_RegFile[27][7]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][7]~q\,
	combout => \Mux115~22_combout\);

-- Location: LABCELL_X62_Y6_N0
\Mux115~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux115~9_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux115~22_combout\)))) # (\R.curInst\(22) & ((!\Mux115~22_combout\ & ((\RegFile[28][7]~q\))) # (\Mux115~22_combout\ & (\RegFile[29][7]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux115~22_combout\)))) # (\R.curInst\(22) & ((!\Mux115~22_combout\ & ((\RegFile[30][7]~q\))) # (\Mux115~22_combout\ & (\RegFile[31][7]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[29][7]~q\,
	datab => \ALT_INV_RegFile[31][7]~q\,
	datac => \ALT_INV_RegFile[30][7]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux115~22_combout\,
	datag => \ALT_INV_RegFile[28][7]~q\,
	combout => \Mux115~9_combout\);

-- Location: LABCELL_X68_Y7_N15
\Mux115~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux115~13_combout\ = ( \Mux115~1_combout\ & ( \Mux115~9_combout\ & ( ((!\R.curInst\(24) & (\Mux115~26_combout\)) # (\R.curInst\(24) & ((\Mux115~5_combout\)))) # (\R.curInst\(23)) ) ) ) # ( !\Mux115~1_combout\ & ( \Mux115~9_combout\ & ( (!\R.curInst\(23) 
-- & ((!\R.curInst\(24) & (\Mux115~26_combout\)) # (\R.curInst\(24) & ((\Mux115~5_combout\))))) # (\R.curInst\(23) & (((\R.curInst\(24))))) ) ) ) # ( \Mux115~1_combout\ & ( !\Mux115~9_combout\ & ( (!\R.curInst\(23) & ((!\R.curInst\(24) & 
-- (\Mux115~26_combout\)) # (\R.curInst\(24) & ((\Mux115~5_combout\))))) # (\R.curInst\(23) & (((!\R.curInst\(24))))) ) ) ) # ( !\Mux115~1_combout\ & ( !\Mux115~9_combout\ & ( (!\R.curInst\(23) & ((!\R.curInst\(24) & (\Mux115~26_combout\)) # (\R.curInst\(24) 
-- & ((\Mux115~5_combout\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010001000001010011101110000101000100010010111110111011101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(23),
	datab => \ALT_INV_Mux115~26_combout\,
	datac => \ALT_INV_Mux115~5_combout\,
	datad => \ALT_INV_R.curInst\(24),
	datae => \ALT_INV_Mux115~1_combout\,
	dataf => \ALT_INV_Mux115~9_combout\,
	combout => \Mux115~13_combout\);

-- Location: LABCELL_X74_Y7_N6
\NxR.aluData2[7]~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[7]~14_combout\ = ( \Mux115~13_combout\ & ( (!\vAluSrc2~1_combout\) # ((\Equal4~1_combout\ & \Mux147~0_combout\)) ) ) # ( !\Mux115~13_combout\ & ( (\vAluSrc2~1_combout\ & (\Equal4~1_combout\ & \Mux147~0_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000011000000000000001111001100110011111100110011001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_vAluSrc2~1_combout\,
	datac => \ALT_INV_Equal4~1_combout\,
	datad => \ALT_INV_Mux147~0_combout\,
	dataf => \ALT_INV_Mux115~13_combout\,
	combout => \NxR.aluData2[7]~14_combout\);

-- Location: FF_X74_Y7_N8
\Add2~25_OTERM723_NEW_REG830\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR.aluData2[7]~14_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Add2~25_OTERM723_OTERM831\);

-- Location: LABCELL_X83_Y5_N24
\vAluRes~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~7_combout\ = ( \vAluRes~7_RESYN1076_BDD1077\ & ( \Add2~29_sumout\ ) ) # ( !\vAluRes~7_RESYN1076_BDD1077\ & ( \Add2~29_sumout\ & ( (\R.aluCalc~q\ & (((\R.aluOp.ALUOpAdd~q\ & \Add1~29_sumout\)) # (\R.aluOp.ALUOpSub~q\))) ) ) ) # ( 
-- \vAluRes~7_RESYN1076_BDD1077\ & ( !\Add2~29_sumout\ ) ) # ( !\vAluRes~7_RESYN1076_BDD1077\ & ( !\Add2~29_sumout\ & ( (\R.aluOp.ALUOpAdd~q\ & (\R.aluCalc~q\ & \Add1~29_sumout\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000101111111111111111100000011000001111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_R.aluCalc~q\,
	datad => \ALT_INV_Add1~29_sumout\,
	datae => \ALT_INV_vAluRes~7_RESYN1076_BDD1077\,
	dataf => \ALT_INV_Add2~29_sumout\,
	combout => \vAluRes~7_combout\);

-- Location: MLABCELL_X84_Y5_N33
\Comb:vJumpAdr[7]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[7]~0_combout\ = ( \Equal4~2_combout\ & ( \Add3~29_sumout\ & ( \vAluRes~7_combout\ ) ) ) # ( !\Equal4~2_combout\ & ( \Add3~29_sumout\ ) ) # ( \Equal4~2_combout\ & ( !\Add3~29_sumout\ & ( \vAluRes~7_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000111111111111111111110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_vAluRes~7_combout\,
	datae => \ALT_INV_Equal4~2_combout\,
	dataf => \ALT_INV_Add3~29_sumout\,
	combout => \Comb:vJumpAdr[7]~0_combout\);

-- Location: FF_X84_Y5_N34
\R.curPC[7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[7]~0_combout\,
	asdata => \Add0~21_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(7));

-- Location: MLABCELL_X78_Y8_N21
\R.regWriteData[8]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.regWriteData[8]~feeder_combout\ = ( \Add0~25_sumout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_Add0~25_sumout\,
	combout => \R.regWriteData[8]~feeder_combout\);

-- Location: LABCELL_X75_Y7_N6
\Selector24~0_RTM0421\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector24~0_RTM0421_combout\ = ( \NxR.aluData2[8]~13_combout\ & ( \R.aluOp.ALUOpAnd_OTERM357\ & ( ((\R.aluOp.ALUOpOr_OTERM353\) # (\Mux246~0_combout\)) # (\R.aluOp.ALUOpXor_OTERM355\) ) ) ) # ( !\NxR.aluData2[8]~13_combout\ & ( 
-- \R.aluOp.ALUOpAnd_OTERM357\ & ( (\Mux246~0_combout\ & ((\R.aluOp.ALUOpOr_OTERM353\) # (\R.aluOp.ALUOpXor_OTERM355\))) ) ) ) # ( \NxR.aluData2[8]~13_combout\ & ( !\R.aluOp.ALUOpAnd_OTERM357\ & ( ((\R.aluOp.ALUOpXor_OTERM355\ & !\Mux246~0_combout\)) # 
-- (\R.aluOp.ALUOpOr_OTERM353\) ) ) ) # ( !\NxR.aluData2[8]~13_combout\ & ( !\R.aluOp.ALUOpAnd_OTERM357\ & ( (\Mux246~0_combout\ & ((\R.aluOp.ALUOpOr_OTERM353\) # (\R.aluOp.ALUOpXor_OTERM355\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100001111010100001111111100000101000011110101111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpXor_OTERM355\,
	datac => \ALT_INV_Mux246~0_combout\,
	datad => \ALT_INV_R.aluOp.ALUOpOr_OTERM353\,
	datae => \ALT_INV_NxR.aluData2[8]~13_combout\,
	dataf => \ALT_INV_R.aluOp.ALUOpAnd_OTERM357\,
	combout => \Selector24~0_RTM0421_combout\);

-- Location: FF_X75_Y7_N7
\Selector24~0_NEW_REG418\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector24~0_RTM0421_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector24~0_OTERM419\);

-- Location: LABCELL_X77_Y8_N30
\Selector24~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector24~1_combout\ = ( \R.aluData1\(31) & ( (!\Selector24~0_OTERM419\ & ((!\R.aluData2\(3)) # (!\Selector31~6_OTERM381\))) ) ) # ( !\R.aluData1\(31) & ( !\Selector24~0_OTERM419\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1100110011001100110011001100110011001100110000001100110011000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Selector24~0_OTERM419\,
	datac => \ALT_INV_R.aluData2\(3),
	datad => \ALT_INV_Selector31~6_OTERM381\,
	dataf => \ALT_INV_R.aluData1\(31),
	combout => \Selector24~1_combout\);

-- Location: MLABCELL_X78_Y8_N18
\Comb:vRegWriteData[8]~1_RESYN1734\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[8]~1_RESYN1734_BDD1735\ = ( \R.memToReg~q\ ) # ( !\R.memToReg~q\ & ( (!\R.aluCalc~q\) # (!\Selector24~1_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111110011111100111111001111110011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_Selector24~1_combout\,
	dataf => \ALT_INV_R.memToReg~q\,
	combout => \Comb:vRegWriteData[8]~1_RESYN1734_BDD1735\);

-- Location: LABCELL_X74_Y8_N45
\ShiftLeft0~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~11_combout\ = ( \R.aluData2\(3) & ( \ShiftLeft0~0_OTERM263\ & ( !\R.aluData2\(2) ) ) ) # ( !\R.aluData2\(3) & ( \ShiftLeft0~0_OTERM263\ & ( (!\R.aluData2\(2) & ((\ShiftLeft0~10_OTERM211\))) # (\R.aluData2\(2) & (\ShiftLeft0~5_OTERM203\)) ) ) ) 
-- # ( !\R.aluData2\(3) & ( !\ShiftLeft0~0_OTERM263\ & ( (!\R.aluData2\(2) & ((\ShiftLeft0~10_OTERM211\))) # (\R.aluData2\(2) & (\ShiftLeft0~5_OTERM203\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111101010101000000000000000000001111010101011111111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~5_OTERM203\,
	datac => \ALT_INV_ShiftLeft0~10_OTERM211\,
	datad => \ALT_INV_R.aluData2\(2),
	datae => \ALT_INV_R.aluData2\(3),
	dataf => \ALT_INV_ShiftLeft0~0_OTERM263\,
	combout => \ShiftLeft0~11_combout\);

-- Location: LABCELL_X74_Y8_N3
\ShiftRight0~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight0~10_combout\ = ( \R.aluData2\(2) & ( (\ShiftRight1~3_OTERM13\ & !\R.aluData2\(3)) ) ) # ( !\R.aluData2\(2) & ( (\ShiftRight1~2_OTERM49\ & !\R.aluData2\(3)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100000000000011110000000001010101000000000101010100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~3_OTERM13\,
	datac => \ALT_INV_ShiftRight1~2_OTERM49\,
	datad => \ALT_INV_R.aluData2\(3),
	dataf => \ALT_INV_R.aluData2\(2),
	combout => \ShiftRight0~10_combout\);

-- Location: LABCELL_X75_Y7_N24
\ShiftRight1~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~7_combout\ = ( \Mux244~0_combout\ & ( \Mux243~0_combout\ & ( ((!\NxR.aluData2[0]~16_combout\ & (\Mux246~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & ((\Mux245~0_combout\)))) # (\NxR.aluData2[1]~17_combout\) ) ) ) # ( !\Mux244~0_combout\ & ( 
-- \Mux243~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((!\NxR.aluData2[0]~16_combout\ & (\Mux246~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & ((\Mux245~0_combout\))))) # (\NxR.aluData2[1]~17_combout\ & (((\NxR.aluData2[0]~16_combout\)))) ) ) ) # ( 
-- \Mux244~0_combout\ & ( !\Mux243~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((!\NxR.aluData2[0]~16_combout\ & (\Mux246~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & ((\Mux245~0_combout\))))) # (\NxR.aluData2[1]~17_combout\ & 
-- (((!\NxR.aluData2[0]~16_combout\)))) ) ) ) # ( !\Mux244~0_combout\ & ( !\Mux243~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((!\NxR.aluData2[0]~16_combout\ & (\Mux246~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & ((\Mux245~0_combout\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100000001001100011100000111110001000011010011110111001101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux246~0_combout\,
	datab => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datac => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datad => \ALT_INV_Mux245~0_combout\,
	datae => \ALT_INV_Mux244~0_combout\,
	dataf => \ALT_INV_Mux243~0_combout\,
	combout => \ShiftRight1~7_combout\);

-- Location: FF_X75_Y7_N25
\ShiftRight1~7_NEW_REG258\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~7_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~7_OTERM259\);

-- Location: LABCELL_X74_Y8_N54
\ShiftRight1~46\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~46_combout\ = ( \R.aluData2\(3) & ( \ShiftRight1~1_OTERM33\ & ( (\R.aluData2\(2)) # (\ShiftRight1~0_OTERM257\) ) ) ) # ( !\R.aluData2\(3) & ( \ShiftRight1~1_OTERM33\ & ( (!\R.aluData2\(2) & (\ShiftRight1~7_OTERM259\)) # (\R.aluData2\(2) & 
-- ((\ShiftRight1~8_OTERM261\))) ) ) ) # ( \R.aluData2\(3) & ( !\ShiftRight1~1_OTERM33\ & ( (\ShiftRight1~0_OTERM257\ & !\R.aluData2\(2)) ) ) ) # ( !\R.aluData2\(3) & ( !\ShiftRight1~1_OTERM33\ & ( (!\R.aluData2\(2) & (\ShiftRight1~7_OTERM259\)) # 
-- (\R.aluData2\(2) & ((\ShiftRight1~8_OTERM261\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011000000111111010100000101000000110000001111110101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~0_OTERM257\,
	datab => \ALT_INV_ShiftRight1~7_OTERM259\,
	datac => \ALT_INV_R.aluData2\(2),
	datad => \ALT_INV_ShiftRight1~8_OTERM261\,
	datae => \ALT_INV_R.aluData2\(3),
	dataf => \ALT_INV_ShiftRight1~1_OTERM33\,
	combout => \ShiftRight1~46_combout\);

-- Location: LABCELL_X75_Y8_N18
\Selector24~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector24~3_combout\ = ( \Selector31~0_OTERM349\ & ( \ShiftRight1~46_combout\ & ( (!\R.aluData2\(4)) # (\ShiftRight0~10_combout\) ) ) ) # ( !\Selector31~0_OTERM349\ & ( \ShiftRight1~46_combout\ & ( (\ShiftLeft0~11_combout\ & (!\R.aluData2\(4) & 
-- \R.aluOp.ALUOpSLL~q\)) ) ) ) # ( \Selector31~0_OTERM349\ & ( !\ShiftRight1~46_combout\ & ( (!\R.aluData2\(4) & (\ShiftLeft0~11_combout\ & ((\R.aluOp.ALUOpSLL~q\)))) # (\R.aluData2\(4) & (((\ShiftRight0~10_combout\)))) ) ) ) # ( !\Selector31~0_OTERM349\ & 
-- ( !\ShiftRight1~46_combout\ & ( (\ShiftLeft0~11_combout\ & (!\R.aluData2\(4) & \R.aluOp.ALUOpSLL~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001000100000000110100011100000000010001001100111111001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~11_combout\,
	datab => \ALT_INV_R.aluData2\(4),
	datac => \ALT_INV_ShiftRight0~10_combout\,
	datad => \ALT_INV_R.aluOp.ALUOpSLL~q\,
	datae => \ALT_INV_Selector31~0_OTERM349\,
	dataf => \ALT_INV_ShiftRight1~46_combout\,
	combout => \Selector24~3_combout\);

-- Location: IOIBUF_X62_Y0_N52
\avm_d_readdata[16]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(16),
	o => \avm_d_readdata[16]~input_o\);

-- Location: LABCELL_X79_Y1_N30
\Comb:vRegWriteData[8]~1_RESYN1730\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[8]~1_RESYN1730_BDD1731\ = ( !\R.curInst\(13) & ( \R.curInst\(12) & ( (\avm_d_readdata[16]~input_o\ & \R.memToReg~q\) ) ) ) # ( \R.curInst\(13) & ( !\R.curInst\(12) & ( (\avm_d_readdata[16]~input_o\ & (\R.memToReg~q\ & 
-- !\R.curInst\(14))) ) ) ) # ( !\R.curInst\(13) & ( !\R.curInst\(12) & ( (\R.memToReg~q\ & (!\R.curInst\(14) & \avm_d_readdata[31]~input_o\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110000000100000001000000010001000100010000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_avm_d_readdata[16]~input_o\,
	datab => \ALT_INV_R.memToReg~q\,
	datac => \ALT_INV_R.curInst\(14),
	datad => \ALT_INV_avm_d_readdata[31]~input_o\,
	datae => \ALT_INV_R.curInst\(13),
	dataf => \ALT_INV_R.curInst\(12),
	combout => \Comb:vRegWriteData[8]~1_RESYN1730_BDD1731\);

-- Location: MLABCELL_X78_Y8_N30
\Comb:vRegWriteData[8]~1_RESYN1732\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[8]~1_RESYN1732_BDD1733\ = ( \R.aluCalc~q\ & ( \Comb:vRegWriteData[8]~1_RESYN1730_BDD1731\ & ( (!\Selector24~1_combout\) # ((\R.aluOp.ALUOpSub~q\) # (\R.memToReg~q\)) ) ) ) # ( !\R.aluCalc~q\ & ( 
-- \Comb:vRegWriteData[8]~1_RESYN1730_BDD1731\ ) ) # ( \R.aluCalc~q\ & ( !\Comb:vRegWriteData[8]~1_RESYN1730_BDD1731\ & ( (!\R.memToReg~q\ & ((!\Selector24~1_combout\) # (\R.aluOp.ALUOpSub~q\))) ) ) ) # ( !\R.aluCalc~q\ & ( 
-- !\Comb:vRegWriteData[8]~1_RESYN1730_BDD1731\ & ( (!\R.memToReg~q\ & \R.aluRes\(8)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011001100100011001000110011111111111111111011111110111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector24~1_combout\,
	datab => \ALT_INV_R.memToReg~q\,
	datac => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datad => \ALT_INV_R.aluRes\(8),
	datae => \ALT_INV_R.aluCalc~q\,
	dataf => \ALT_INV_Comb:vRegWriteData[8]~1_RESYN1730_BDD1731\,
	combout => \Comb:vRegWriteData[8]~1_RESYN1732_BDD1733\);

-- Location: MLABCELL_X78_Y8_N54
\Comb:vRegWriteData[8]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[8]~1_combout\ = ( \Add2~33_sumout\ & ( \Comb:vRegWriteData[8]~1_RESYN1732_BDD1733\ ) ) # ( !\Add2~33_sumout\ & ( \Comb:vRegWriteData[8]~1_RESYN1732_BDD1733\ & ( (((\R.aluOp.ALUOpAdd~q\ & \Add1~33_sumout\)) # (\Selector24~3_combout\)) # 
-- (\Comb:vRegWriteData[8]~1_RESYN1734_BDD1735\) ) ) ) # ( \Add2~33_sumout\ & ( !\Comb:vRegWriteData[8]~1_RESYN1732_BDD1733\ & ( (!\Comb:vRegWriteData[8]~1_RESYN1734_BDD1735\ & (((\R.aluOp.ALUOpAdd~q\ & \Add1~33_sumout\)) # (\Selector24~3_combout\))) ) ) ) # 
-- ( !\Add2~33_sumout\ & ( !\Comb:vRegWriteData[8]~1_RESYN1732_BDD1733\ & ( (!\Comb:vRegWriteData[8]~1_RESYN1734_BDD1735\ & (((\R.aluOp.ALUOpAdd~q\ & \Add1~33_sumout\)) # (\Selector24~3_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101000101010000010100010101001011111011111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Comb:vRegWriteData[8]~1_RESYN1734_BDD1735\,
	datab => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datac => \ALT_INV_Selector24~3_combout\,
	datad => \ALT_INV_Add1~33_sumout\,
	datae => \ALT_INV_Add2~33_sumout\,
	dataf => \ALT_INV_Comb:vRegWriteData[8]~1_RESYN1732_BDD1733\,
	combout => \Comb:vRegWriteData[8]~1_combout\);

-- Location: FF_X78_Y8_N23
\R.regWriteData[8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \R.regWriteData[8]~feeder_combout\,
	asdata => \Comb:vRegWriteData[8]~1_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(8));

-- Location: FF_X67_Y7_N32
\RegFile[3][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(8),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][8]~q\);

-- Location: FF_X65_Y7_N56
\RegFile[2][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(8),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][8]~q\);

-- Location: LABCELL_X55_Y7_N0
\RegFile[5][8]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[5][8]~feeder_combout\ = ( \R.regWriteData\(8) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(8),
	combout => \RegFile[5][8]~feeder_combout\);

-- Location: FF_X55_Y7_N1
\RegFile[5][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[5][8]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][8]~q\);

-- Location: LABCELL_X67_Y7_N36
\RegFile[6][8]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[6][8]~feeder_combout\ = ( \R.regWriteData\(8) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(8),
	combout => \RegFile[6][8]~feeder_combout\);

-- Location: FF_X67_Y7_N37
\RegFile[6][8]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[6][8]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][8]~DUPLICATE_q\);

-- Location: FF_X67_Y5_N19
\RegFile[4][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(8),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][8]~q\);

-- Location: FF_X67_Y7_N44
\RegFile[7][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(8),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][8]~q\);

-- Location: MLABCELL_X65_Y7_N39
\Mux114~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux114~0_combout\ = ( \RegFile[7][8]~q\ & ( \R.curInst\(21) & ( (\R.curInst\(20)) # (\RegFile[6][8]~DUPLICATE_q\) ) ) ) # ( !\RegFile[7][8]~q\ & ( \R.curInst\(21) & ( (\RegFile[6][8]~DUPLICATE_q\ & !\R.curInst\(20)) ) ) ) # ( \RegFile[7][8]~q\ & ( 
-- !\R.curInst\(21) & ( (!\R.curInst\(20) & ((\RegFile[4][8]~q\))) # (\R.curInst\(20) & (\RegFile[5][8]~q\)) ) ) ) # ( !\RegFile[7][8]~q\ & ( !\R.curInst\(21) & ( (!\R.curInst\(20) & ((\RegFile[4][8]~q\))) # (\R.curInst\(20) & (\RegFile[5][8]~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111101010101000011110101010100110011000000000011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[5][8]~q\,
	datab => \ALT_INV_RegFile[6][8]~DUPLICATE_q\,
	datac => \ALT_INV_RegFile[4][8]~q\,
	datad => \ALT_INV_R.curInst\(20),
	datae => \ALT_INV_RegFile[7][8]~q\,
	dataf => \ALT_INV_R.curInst\(21),
	combout => \Mux114~0_combout\);

-- Location: MLABCELL_X59_Y7_N12
\RegFile[1][8]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[1][8]~feeder_combout\ = ( \R.regWriteData\(8) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(8),
	combout => \RegFile[1][8]~feeder_combout\);

-- Location: FF_X59_Y7_N13
\RegFile[1][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[1][8]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][8]~q\);

-- Location: MLABCELL_X65_Y7_N54
\Mux114~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux114~26_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (\R.curInst\(20) & (\RegFile[1][8]~q\))) # (\R.curInst\(22) & (((\Mux114~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (((\RegFile[2][8]~q\)))) # 
-- (\R.curInst\(20) & (\RegFile[3][8]~q\)))) # (\R.curInst\(22) & ((((\Mux114~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000000000111010000000000000011111111110001110111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][8]~q\,
	datab => \ALT_INV_R.curInst\(20),
	datac => \ALT_INV_RegFile[2][8]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux114~0_combout\,
	datag => \ALT_INV_RegFile[1][8]~q\,
	combout => \Mux114~26_combout\);

-- Location: FF_X66_Y7_N50
\RegFile[13][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(8),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][8]~q\);

-- Location: FF_X62_Y9_N55
\RegFile[14][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(8),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][8]~q\);

-- Location: FF_X66_Y7_N8
\RegFile[15][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(8),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][8]~q\);

-- Location: FF_X65_Y3_N2
\RegFile[9][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(8),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][8]~q\);

-- Location: MLABCELL_X65_Y3_N6
\RegFile[11][8]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[11][8]~feeder_combout\ = ( \R.regWriteData\(8) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(8),
	combout => \RegFile[11][8]~feeder_combout\);

-- Location: FF_X65_Y3_N8
\RegFile[11][8]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[11][8]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][8]~DUPLICATE_q\);

-- Location: MLABCELL_X65_Y3_N48
\RegFile[10][8]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[10][8]~feeder_combout\ = ( \R.regWriteData\(8) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(8),
	combout => \RegFile[10][8]~feeder_combout\);

-- Location: FF_X65_Y3_N49
\RegFile[10][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[10][8]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][8]~q\);

-- Location: LABCELL_X55_Y5_N39
\RegFile[8][8]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[8][8]~feeder_combout\ = ( \R.regWriteData\(8) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(8),
	combout => \RegFile[8][8]~feeder_combout\);

-- Location: FF_X55_Y5_N40
\RegFile[8][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[8][8]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][8]~q\);

-- Location: MLABCELL_X65_Y3_N0
\Mux114~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux114~14_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[8][8]~q\))) # (\R.curInst\(20) & (\RegFile[9][8]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[10][8]~q\))) # (\R.curInst\(20) & (\RegFile[11][8]~DUPLICATE_q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][8]~q\,
	datab => \ALT_INV_RegFile[11][8]~DUPLICATE_q\,
	datac => \ALT_INV_RegFile[10][8]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][8]~q\,
	combout => \Mux114~14_combout\);

-- Location: LABCELL_X66_Y7_N36
\RegFile[12][8]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[12][8]~feeder_combout\ = ( \R.regWriteData\(8) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(8),
	combout => \RegFile[12][8]~feeder_combout\);

-- Location: FF_X66_Y7_N38
\RegFile[12][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[12][8]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][8]~q\);

-- Location: LABCELL_X66_Y7_N48
\Mux114~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux114~1_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux114~14_combout\))))) # (\R.curInst\(22) & (((!\Mux114~14_combout\ & ((\RegFile[12][8]~q\))) # (\Mux114~14_combout\ & (\RegFile[13][8]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux114~14_combout\)))) # (\R.curInst\(22) & ((!\Mux114~14_combout\ & (\RegFile[14][8]~q\)) # (\Mux114~14_combout\ & ((\RegFile[15][8]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][8]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[14][8]~q\,
	datad => \ALT_INV_RegFile[15][8]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux114~14_combout\,
	datag => \ALT_INV_RegFile[12][8]~q\,
	combout => \Mux114~1_combout\);

-- Location: FF_X65_Y8_N2
\RegFile[21][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(8),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][8]~q\);

-- Location: FF_X64_Y4_N38
\RegFile[23][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(8),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][8]~q\);

-- Location: LABCELL_X64_Y4_N3
\RegFile[22][8]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[22][8]~feeder_combout\ = ( \R.regWriteData\(8) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(8),
	combout => \RegFile[22][8]~feeder_combout\);

-- Location: FF_X64_Y4_N5
\RegFile[22][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[22][8]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][8]~q\);

-- Location: FF_X65_Y8_N44
\RegFile[17][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(8),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][8]~q\);

-- Location: FF_X64_Y4_N50
\RegFile[19][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(8),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][8]~q\);

-- Location: LABCELL_X64_Y10_N6
\RegFile[18][8]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[18][8]~feeder_combout\ = ( \R.regWriteData\(8) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(8),
	combout => \RegFile[18][8]~feeder_combout\);

-- Location: FF_X64_Y10_N7
\RegFile[18][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][8]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][8]~q\);

-- Location: LABCELL_X55_Y7_N27
\RegFile[16][8]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[16][8]~feeder_combout\ = ( \R.regWriteData\(8) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(8),
	combout => \RegFile[16][8]~feeder_combout\);

-- Location: FF_X55_Y7_N28
\RegFile[16][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[16][8]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][8]~q\);

-- Location: MLABCELL_X65_Y8_N42
\Mux114~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux114~18_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[16][8]~q\))) # (\R.curInst\(20) & (\RegFile[17][8]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[18][8]~q\))) # (\R.curInst\(20) & (\RegFile[19][8]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[17][8]~q\,
	datab => \ALT_INV_RegFile[19][8]~q\,
	datac => \ALT_INV_RegFile[18][8]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][8]~q\,
	combout => \Mux114~18_combout\);

-- Location: LABCELL_X64_Y10_N54
\RegFile[20][8]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[20][8]~feeder_combout\ = ( \R.regWriteData\(8) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(8),
	combout => \RegFile[20][8]~feeder_combout\);

-- Location: FF_X64_Y10_N55
\RegFile[20][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[20][8]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][8]~q\);

-- Location: MLABCELL_X65_Y8_N0
\Mux114~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux114~5_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux114~18_combout\)))) # (\R.curInst\(22) & ((!\Mux114~18_combout\ & ((\RegFile[20][8]~q\))) # (\Mux114~18_combout\ & (\RegFile[21][8]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux114~18_combout\)))) # (\R.curInst\(22) & ((!\Mux114~18_combout\ & ((\RegFile[22][8]~q\))) # (\Mux114~18_combout\ & (\RegFile[23][8]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][8]~q\,
	datab => \ALT_INV_RegFile[23][8]~q\,
	datac => \ALT_INV_RegFile[22][8]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux114~18_combout\,
	datag => \ALT_INV_RegFile[20][8]~q\,
	combout => \Mux114~5_combout\);

-- Location: FF_X60_Y7_N53
\RegFile[29][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(8),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][8]~q\);

-- Location: LABCELL_X60_Y7_N12
\RegFile[31][8]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[31][8]~feeder_combout\ = ( \R.regWriteData\(8) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(8),
	combout => \RegFile[31][8]~feeder_combout\);

-- Location: FF_X60_Y7_N14
\RegFile[31][8]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[31][8]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][8]~DUPLICATE_q\);

-- Location: LABCELL_X55_Y7_N6
\RegFile[30][8]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[30][8]~feeder_combout\ = ( \R.regWriteData\(8) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(8),
	combout => \RegFile[30][8]~feeder_combout\);

-- Location: FF_X55_Y7_N7
\RegFile[30][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[30][8]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][8]~q\);

-- Location: FF_X61_Y3_N32
\RegFile[27][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(8),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][8]~q\);

-- Location: FF_X57_Y6_N58
\RegFile[26][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(8),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][8]~q\);

-- Location: LABCELL_X61_Y3_N54
\RegFile[25][8]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[25][8]~feeder_combout\ = ( \R.regWriteData\(8) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(8),
	combout => \RegFile[25][8]~feeder_combout\);

-- Location: FF_X61_Y3_N55
\RegFile[25][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[25][8]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][8]~q\);

-- Location: LABCELL_X56_Y3_N33
\RegFile[24][8]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[24][8]~feeder_combout\ = ( \R.regWriteData\(8) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(8),
	combout => \RegFile[24][8]~feeder_combout\);

-- Location: FF_X56_Y3_N34
\RegFile[24][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[24][8]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][8]~q\);

-- Location: LABCELL_X60_Y7_N39
\Mux114~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux114~22_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & (\RegFile[24][8]~q\)) # (\R.curInst\(20) & ((\RegFile[25][8]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & ((\RegFile[26][8]~q\))) # (\R.curInst\(20) & (\RegFile[27][8]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110000110011111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[27][8]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[26][8]~q\,
	datad => \ALT_INV_RegFile[25][8]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][8]~q\,
	combout => \Mux114~22_combout\);

-- Location: MLABCELL_X65_Y9_N15
\RegFile[28][8]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[28][8]~feeder_combout\ = ( \R.regWriteData\(8) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(8),
	combout => \RegFile[28][8]~feeder_combout\);

-- Location: FF_X65_Y9_N16
\RegFile[28][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[28][8]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][8]~q\);

-- Location: LABCELL_X60_Y7_N51
\Mux114~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux114~9_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux114~22_combout\)))) # (\R.curInst\(22) & ((!\Mux114~22_combout\ & ((\RegFile[28][8]~q\))) # (\Mux114~22_combout\ & (\RegFile[29][8]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux114~22_combout\)))) # (\R.curInst\(22) & ((!\Mux114~22_combout\ & ((\RegFile[30][8]~q\))) # (\Mux114~22_combout\ & (\RegFile[31][8]~DUPLICATE_q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[29][8]~q\,
	datab => \ALT_INV_RegFile[31][8]~DUPLICATE_q\,
	datac => \ALT_INV_RegFile[30][8]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux114~22_combout\,
	datag => \ALT_INV_RegFile[28][8]~q\,
	combout => \Mux114~9_combout\);

-- Location: MLABCELL_X65_Y7_N42
\Mux114~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux114~13_combout\ = ( \Mux114~5_combout\ & ( \Mux114~9_combout\ & ( ((!\R.curInst\(23) & (\Mux114~26_combout\)) # (\R.curInst\(23) & ((\Mux114~1_combout\)))) # (\R.curInst\(24)) ) ) ) # ( !\Mux114~5_combout\ & ( \Mux114~9_combout\ & ( (!\R.curInst\(23) 
-- & (\Mux114~26_combout\ & (!\R.curInst\(24)))) # (\R.curInst\(23) & (((\Mux114~1_combout\) # (\R.curInst\(24))))) ) ) ) # ( \Mux114~5_combout\ & ( !\Mux114~9_combout\ & ( (!\R.curInst\(23) & (((\R.curInst\(24))) # (\Mux114~26_combout\))) # (\R.curInst\(23) 
-- & (((!\R.curInst\(24) & \Mux114~1_combout\)))) ) ) ) # ( !\Mux114~5_combout\ & ( !\Mux114~9_combout\ & ( (!\R.curInst\(24) & ((!\R.curInst\(23) & (\Mux114~26_combout\)) # (\R.curInst\(23) & ((\Mux114~1_combout\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010000001110000001010100111101000100101011101010010111101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(23),
	datab => \ALT_INV_Mux114~26_combout\,
	datac => \ALT_INV_R.curInst\(24),
	datad => \ALT_INV_Mux114~1_combout\,
	datae => \ALT_INV_Mux114~5_combout\,
	dataf => \ALT_INV_Mux114~9_combout\,
	combout => \Mux114~13_combout\);

-- Location: LABCELL_X74_Y7_N27
\NxR.aluData2[8]~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[8]~13_combout\ = ( \Mux114~13_combout\ & ( (!\vAluSrc2~1_combout\) # ((\Equal4~1_combout\ & \Mux146~0_combout\)) ) ) # ( !\Mux114~13_combout\ & ( (\Equal4~1_combout\ & (\vAluSrc2~1_combout\ & \Mux146~0_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000101000000000000010111110000111101011111000011110101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Equal4~1_combout\,
	datac => \ALT_INV_vAluSrc2~1_combout\,
	datad => \ALT_INV_Mux146~0_combout\,
	dataf => \ALT_INV_Mux114~13_combout\,
	combout => \NxR.aluData2[8]~13_combout\);

-- Location: FF_X74_Y7_N16
\Add2~33_OTERM719_NEW_REG826\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \NxR.aluData2[8]~13_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Add2~33_OTERM719_OTERM827\);

-- Location: LABCELL_X79_Y8_N0
\Selector24~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector24~4_combout\ = ( \R.aluOp.ALUOpAdd~q\ & ( \Add2~33_sumout\ & ( (((!\Selector24~1_combout\) # (\Selector24~3_combout\)) # (\Add1~33_sumout\)) # (\R.aluOp.ALUOpSub~q\) ) ) ) # ( !\R.aluOp.ALUOpAdd~q\ & ( \Add2~33_sumout\ & ( 
-- ((!\Selector24~1_combout\) # (\Selector24~3_combout\)) # (\R.aluOp.ALUOpSub~q\) ) ) ) # ( \R.aluOp.ALUOpAdd~q\ & ( !\Add2~33_sumout\ & ( ((!\Selector24~1_combout\) # (\Selector24~3_combout\)) # (\Add1~33_sumout\) ) ) ) # ( !\R.aluOp.ALUOpAdd~q\ & ( 
-- !\Add2~33_sumout\ & ( (!\Selector24~1_combout\) # (\Selector24~3_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111000011111111111100111111111111110101111111111111011111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datab => \ALT_INV_Add1~33_sumout\,
	datac => \ALT_INV_Selector24~1_combout\,
	datad => \ALT_INV_Selector24~3_combout\,
	datae => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	dataf => \ALT_INV_Add2~33_sumout\,
	combout => \Selector24~4_combout\);

-- Location: FF_X79_Y8_N1
\R.aluRes[8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector24~4_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(8));

-- Location: LABCELL_X80_Y8_N24
\vAluRes~31\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~31_combout\ = ( \Selector24~3_combout\ & ( (!\R.aluRes\(8) & !\R.aluCalc~q\) ) ) # ( !\Selector24~3_combout\ & ( (!\R.aluCalc~q\ & (!\R.aluRes\(8))) # (\R.aluCalc~q\ & ((\Selector24~1_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010101000001111101010100000111110101010000000001010101000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluRes\(8),
	datac => \ALT_INV_Selector24~1_combout\,
	datad => \ALT_INV_R.aluCalc~q\,
	dataf => \ALT_INV_Selector24~3_combout\,
	combout => \vAluRes~31_combout\);

-- Location: LABCELL_X79_Y8_N54
\vAluRes~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~8_combout\ = ( \Add1~33_sumout\ & ( \Add2~33_sumout\ & ( (!\vAluRes~31_combout\) # ((\R.aluCalc~q\ & ((\R.aluOp.ALUOpAdd~q\) # (\R.aluOp.ALUOpSub~q\)))) ) ) ) # ( !\Add1~33_sumout\ & ( \Add2~33_sumout\ & ( (!\vAluRes~31_combout\) # 
-- ((\R.aluOp.ALUOpSub~q\ & \R.aluCalc~q\)) ) ) ) # ( \Add1~33_sumout\ & ( !\Add2~33_sumout\ & ( (!\vAluRes~31_combout\) # ((\R.aluCalc~q\ & \R.aluOp.ALUOpAdd~q\)) ) ) ) # ( !\Add1~33_sumout\ & ( !\Add2~33_sumout\ & ( !\vAluRes~31_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111100000000111111110000001111111111000100011111111100010011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_vAluRes~31_combout\,
	datae => \ALT_INV_Add1~33_sumout\,
	dataf => \ALT_INV_Add2~33_sumout\,
	combout => \vAluRes~8_combout\);

-- Location: MLABCELL_X78_Y8_N42
\Comb:vJumpAdr[8]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[8]~0_combout\ = ( \Equal4~2_combout\ & ( \Add3~33_sumout\ & ( \vAluRes~8_combout\ ) ) ) # ( !\Equal4~2_combout\ & ( \Add3~33_sumout\ ) ) # ( \Equal4~2_combout\ & ( !\Add3~33_sumout\ & ( \vAluRes~8_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000001100110011001111111111111111110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_vAluRes~8_combout\,
	datae => \ALT_INV_Equal4~2_combout\,
	dataf => \ALT_INV_Add3~33_sumout\,
	combout => \Comb:vJumpAdr[8]~0_combout\);

-- Location: FF_X78_Y8_N43
\R.curPC[8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[8]~0_combout\,
	asdata => \Add0~25_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(8));

-- Location: FF_X60_Y7_N13
\RegFile[31][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[31][8]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][8]~q\);

-- Location: LABCELL_X61_Y3_N30
\Mux82~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux82~22_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & (\RegFile[24][8]~q\)) # (\R.curInst\(15) & ((\RegFile[25][8]~q\)))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & ((\RegFile[26][8]~q\))) # (\R.curInst\(15) & (\RegFile[27][8]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001010101111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[27][8]~q\,
	datac => \ALT_INV_RegFile[26][8]~q\,
	datad => \ALT_INV_RegFile[25][8]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][8]~q\,
	combout => \Mux82~22_combout\);

-- Location: LABCELL_X73_Y7_N12
\Mux82~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux82~9_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux82~22_combout\)))) # (\R.curInst\(17) & ((!\Mux82~22_combout\ & ((\RegFile[28][8]~q\))) # (\Mux82~22_combout\ & (\RegFile[29][8]~q\))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) 
-- & (((\Mux82~22_combout\)))) # (\R.curInst\(17) & ((!\Mux82~22_combout\ & ((\RegFile[30][8]~q\))) # (\Mux82~22_combout\ & (\RegFile[31][8]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[29][8]~q\,
	datab => \ALT_INV_RegFile[31][8]~q\,
	datac => \ALT_INV_RegFile[30][8]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux82~22_combout\,
	datag => \ALT_INV_RegFile[28][8]~q\,
	combout => \Mux82~9_combout\);

-- Location: FF_X67_Y7_N38
\RegFile[6][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[6][8]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][8]~q\);

-- Location: LABCELL_X67_Y7_N42
\Mux82~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux82~0_combout\ = ( \RegFile[7][8]~q\ & ( \R.curInst\(15) & ( (\RegFile[5][8]~q\) # (\R.curInst\(16)) ) ) ) # ( !\RegFile[7][8]~q\ & ( \R.curInst\(15) & ( (!\R.curInst\(16) & \RegFile[5][8]~q\) ) ) ) # ( \RegFile[7][8]~q\ & ( !\R.curInst\(15) & ( 
-- (!\R.curInst\(16) & (\RegFile[4][8]~q\)) # (\R.curInst\(16) & ((\RegFile[6][8]~q\))) ) ) ) # ( !\RegFile[7][8]~q\ & ( !\R.curInst\(15) & ( (!\R.curInst\(16) & (\RegFile[4][8]~q\)) # (\R.curInst\(16) & ((\RegFile[6][8]~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100011101000111010001110100011100000000110011000011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[4][8]~q\,
	datab => \ALT_INV_R.curInst\(16),
	datac => \ALT_INV_RegFile[6][8]~q\,
	datad => \ALT_INV_RegFile[5][8]~q\,
	datae => \ALT_INV_RegFile[7][8]~q\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux82~0_combout\);

-- Location: LABCELL_X67_Y7_N30
\Mux82~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux82~26_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (\R.curInst\(15) & (\RegFile[1][8]~q\))) # (\R.curInst\(17) & (((\Mux82~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & ((!\R.curInst\(15) & (((\RegFile[2][8]~q\)))) # 
-- (\R.curInst\(15) & (\RegFile[3][8]~q\)))) # (\R.curInst\(17) & ((((\Mux82~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000000000110110000000000000101111111110001101111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(15),
	datab => \ALT_INV_RegFile[3][8]~q\,
	datac => \ALT_INV_RegFile[2][8]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux82~0_combout\,
	datag => \ALT_INV_RegFile[1][8]~q\,
	combout => \Mux82~26_combout\);

-- Location: FF_X65_Y3_N7
\RegFile[11][8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[11][8]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][8]~q\);

-- Location: MLABCELL_X65_Y7_N18
\Mux82~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux82~14_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[8][8]~q\))) # (\R.curInst\(15) & (\RegFile[9][8]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[10][8]~q\))) # (\R.curInst\(15) & (\RegFile[11][8]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[11][8]~q\,
	datab => \ALT_INV_RegFile[9][8]~q\,
	datac => \ALT_INV_RegFile[10][8]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][8]~q\,
	combout => \Mux82~14_combout\);

-- Location: LABCELL_X66_Y7_N6
\Mux82~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux82~1_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux82~14_combout\))))) # (\R.curInst\(17) & (((!\Mux82~14_combout\ & ((\RegFile[12][8]~q\))) # (\Mux82~14_combout\ & (\RegFile[13][8]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux82~14_combout\)))) # (\R.curInst\(17) & ((!\Mux82~14_combout\ & (\RegFile[14][8]~q\)) # (\Mux82~14_combout\ & ((\RegFile[15][8]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][8]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[14][8]~q\,
	datad => \ALT_INV_RegFile[15][8]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux82~14_combout\,
	datag => \ALT_INV_RegFile[12][8]~q\,
	combout => \Mux82~1_combout\);

-- Location: FF_X64_Y10_N8
\RegFile[18][8]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][8]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][8]~DUPLICATE_q\);

-- Location: LABCELL_X64_Y4_N48
\Mux82~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux82~18_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[16][8]~q\))) # (\R.curInst\(15) & (\RegFile[17][8]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[18][8]~DUPLICATE_q\))) # (\R.curInst\(15) & (\RegFile[19][8]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[19][8]~q\,
	datab => \ALT_INV_RegFile[17][8]~q\,
	datac => \ALT_INV_RegFile[18][8]~DUPLICATE_q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][8]~q\,
	combout => \Mux82~18_combout\);

-- Location: LABCELL_X64_Y4_N36
\Mux82~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux82~5_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux82~18_combout\)))) # (\R.curInst\(17) & ((!\Mux82~18_combout\ & ((\RegFile[20][8]~q\))) # (\Mux82~18_combout\ & (\RegFile[21][8]~q\))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) 
-- & (((\Mux82~18_combout\)))) # (\R.curInst\(17) & ((!\Mux82~18_combout\ & ((\RegFile[22][8]~q\))) # (\Mux82~18_combout\ & (\RegFile[23][8]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[23][8]~q\,
	datab => \ALT_INV_RegFile[21][8]~q\,
	datac => \ALT_INV_RegFile[22][8]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux82~18_combout\,
	datag => \ALT_INV_RegFile[20][8]~q\,
	combout => \Mux82~5_combout\);

-- Location: LABCELL_X73_Y7_N54
\Mux82~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux82~13_combout\ = ( \Mux82~1_combout\ & ( \Mux82~5_combout\ & ( (!\R.curInst\(19) & (((\Mux82~26_combout\) # (\R.curInst\(18))))) # (\R.curInst\(19) & (((!\R.curInst\(18))) # (\Mux82~9_combout\))) ) ) ) # ( !\Mux82~1_combout\ & ( \Mux82~5_combout\ & ( 
-- (!\R.curInst\(19) & (((!\R.curInst\(18) & \Mux82~26_combout\)))) # (\R.curInst\(19) & (((!\R.curInst\(18))) # (\Mux82~9_combout\))) ) ) ) # ( \Mux82~1_combout\ & ( !\Mux82~5_combout\ & ( (!\R.curInst\(19) & (((\Mux82~26_combout\) # (\R.curInst\(18))))) # 
-- (\R.curInst\(19) & (\Mux82~9_combout\ & (\R.curInst\(18)))) ) ) ) # ( !\Mux82~1_combout\ & ( !\Mux82~5_combout\ & ( (!\R.curInst\(19) & (((!\R.curInst\(18) & \Mux82~26_combout\)))) # (\R.curInst\(19) & (\Mux82~9_combout\ & (\R.curInst\(18)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000110100001000010111010101101010001111100010101101111111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(19),
	datab => \ALT_INV_Mux82~9_combout\,
	datac => \ALT_INV_R.curInst\(18),
	datad => \ALT_INV_Mux82~26_combout\,
	datae => \ALT_INV_Mux82~1_combout\,
	dataf => \ALT_INV_Mux82~5_combout\,
	combout => \Mux82~13_combout\);

-- Location: LABCELL_X74_Y7_N54
\Mux246~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux246~0_combout\ = ( \Mux82~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC\(8)))) ) ) # ( !\Mux82~13_combout\ & ( (!\vAluSrc1~1_combout\ & (\vAluSrc1~2_combout\ & \R.curPC\(8))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001000000010000000100000001010001010100010101000101010001010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluSrc1~1_combout\,
	datab => \ALT_INV_vAluSrc1~2_combout\,
	datac => \ALT_INV_R.curPC\(8),
	dataf => \ALT_INV_Mux82~13_combout\,
	combout => \Mux246~0_combout\);

-- Location: LABCELL_X75_Y7_N54
\ShiftLeft0~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~14_combout\ = ( \Mux244~0_combout\ & ( \Mux243~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\) # ((!\NxR.aluData2[0]~16_combout\ & ((\Mux245~0_combout\))) # (\NxR.aluData2[0]~16_combout\ & (\Mux246~0_combout\))) ) ) ) # ( !\Mux244~0_combout\ & 
-- ( \Mux243~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((!\NxR.aluData2[0]~16_combout\)))) # (\NxR.aluData2[1]~17_combout\ & ((!\NxR.aluData2[0]~16_combout\ & ((\Mux245~0_combout\))) # (\NxR.aluData2[0]~16_combout\ & (\Mux246~0_combout\)))) ) ) ) # ( 
-- \Mux244~0_combout\ & ( !\Mux243~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((\NxR.aluData2[0]~16_combout\)))) # (\NxR.aluData2[1]~17_combout\ & ((!\NxR.aluData2[0]~16_combout\ & ((\Mux245~0_combout\))) # (\NxR.aluData2[0]~16_combout\ & 
-- (\Mux246~0_combout\)))) ) ) ) # ( !\Mux244~0_combout\ & ( !\Mux243~0_combout\ & ( (\NxR.aluData2[1]~17_combout\ & ((!\NxR.aluData2[0]~16_combout\ & ((\Mux245~0_combout\))) # (\NxR.aluData2[0]~16_combout\ & (\Mux246~0_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000100110001000011010011110111000001111100011100110111111101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux246~0_combout\,
	datab => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datac => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datad => \ALT_INV_Mux245~0_combout\,
	datae => \ALT_INV_Mux244~0_combout\,
	dataf => \ALT_INV_Mux243~0_combout\,
	combout => \ShiftLeft0~14_combout\);

-- Location: FF_X75_Y7_N55
\ShiftLeft0~14_NEW_REG752\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~14_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~14_OTERM753\);

-- Location: LABCELL_X77_Y8_N42
\ShiftLeft0~31\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~31_combout\ = ( \ShiftLeft0~9_OTERM461\ & ( \ShiftLeft0~22_OTERM737\ & ( ((!\R.aluData2\(3) & ((\ShiftLeft0~30_OTERM601\))) # (\R.aluData2\(3) & (\ShiftLeft0~14_OTERM753\))) # (\R.aluData2\(2)) ) ) ) # ( !\ShiftLeft0~9_OTERM461\ & ( 
-- \ShiftLeft0~22_OTERM737\ & ( (!\R.aluData2\(3) & (((\ShiftLeft0~30_OTERM601\)) # (\R.aluData2\(2)))) # (\R.aluData2\(3) & (!\R.aluData2\(2) & (\ShiftLeft0~14_OTERM753\))) ) ) ) # ( \ShiftLeft0~9_OTERM461\ & ( !\ShiftLeft0~22_OTERM737\ & ( 
-- (!\R.aluData2\(3) & (!\R.aluData2\(2) & ((\ShiftLeft0~30_OTERM601\)))) # (\R.aluData2\(3) & (((\ShiftLeft0~14_OTERM753\)) # (\R.aluData2\(2)))) ) ) ) # ( !\ShiftLeft0~9_OTERM461\ & ( !\ShiftLeft0~22_OTERM737\ & ( (!\R.aluData2\(2) & ((!\R.aluData2\(3) & 
-- ((\ShiftLeft0~30_OTERM601\))) # (\R.aluData2\(3) & (\ShiftLeft0~14_OTERM753\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010010001100000101011001110100100110101011100011011110111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(3),
	datab => \ALT_INV_R.aluData2\(2),
	datac => \ALT_INV_ShiftLeft0~14_OTERM753\,
	datad => \ALT_INV_ShiftLeft0~30_OTERM601\,
	datae => \ALT_INV_ShiftLeft0~9_OTERM461\,
	dataf => \ALT_INV_ShiftLeft0~22_OTERM737\,
	combout => \ShiftLeft0~31_combout\);

-- Location: LABCELL_X77_Y7_N3
\ShiftRight1~33\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~33_combout\ = ( \R.aluData2\(3) & ( \R.aluData1\(31) & ( (\ShiftRight1~32_OTERM21\) # (\R.aluData2\(2)) ) ) ) # ( !\R.aluData2\(3) & ( \R.aluData1\(31) & ( (!\R.aluData2\(2) & ((\ShiftRight1~30_OTERM39\))) # (\R.aluData2\(2) & 
-- (\ShiftRight1~31_OTERM45\)) ) ) ) # ( \R.aluData2\(3) & ( !\R.aluData1\(31) & ( (!\R.aluData2\(2) & \ShiftRight1~32_OTERM21\) ) ) ) # ( !\R.aluData2\(3) & ( !\R.aluData1\(31) & ( (!\R.aluData2\(2) & ((\ShiftRight1~30_OTERM39\))) # (\R.aluData2\(2) & 
-- (\ShiftRight1~31_OTERM45\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000111011101000011000000110000010001110111010011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~31_OTERM45\,
	datab => \ALT_INV_R.aluData2\(2),
	datac => \ALT_INV_ShiftRight1~32_OTERM21\,
	datad => \ALT_INV_ShiftRight1~30_OTERM39\,
	datae => \ALT_INV_R.aluData2\(3),
	dataf => \ALT_INV_R.aluData1\(31),
	combout => \ShiftRight1~33_combout\);

-- Location: LABCELL_X77_Y7_N0
\ShiftRight0~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight0~5_combout\ = ( \R.aluData2\(3) & ( \ShiftRight0~4_OTERM31\ & ( (\ShiftRight1~32_OTERM21\) # (\R.aluData2\(2)) ) ) ) # ( !\R.aluData2\(3) & ( \ShiftRight0~4_OTERM31\ & ( (!\R.aluData2\(2) & ((\ShiftRight1~30_OTERM39\))) # (\R.aluData2\(2) & 
-- (\ShiftRight1~31_OTERM45\)) ) ) ) # ( \R.aluData2\(3) & ( !\ShiftRight0~4_OTERM31\ & ( (!\R.aluData2\(2) & \ShiftRight1~32_OTERM21\) ) ) ) # ( !\R.aluData2\(3) & ( !\ShiftRight0~4_OTERM31\ & ( (!\R.aluData2\(2) & ((\ShiftRight1~30_OTERM39\))) # 
-- (\R.aluData2\(2) & (\ShiftRight1~31_OTERM45\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001110100011101000000001100110000011101000111010011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~31_OTERM45\,
	datab => \ALT_INV_R.aluData2\(2),
	datac => \ALT_INV_ShiftRight1~30_OTERM39\,
	datad => \ALT_INV_ShiftRight1~32_OTERM21\,
	datae => \ALT_INV_R.aluData2\(3),
	dataf => \ALT_INV_ShiftRight0~4_OTERM31\,
	combout => \ShiftRight0~5_combout\);

-- Location: MLABCELL_X82_Y5_N27
\Selector13~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector13~0_combout\ = ( \R.aluOp.ALUOpSRA~q\ & ( \ShiftRight0~5_combout\ & ( (!\R.aluOp.ALUOpSRL~q\ & (!\ShiftRight1~33_combout\ & ((!\ShiftLeft0~31_combout\) # (!\R.aluOp.ALUOpSLL~q\)))) ) ) ) # ( !\R.aluOp.ALUOpSRA~q\ & ( \ShiftRight0~5_combout\ & ( 
-- (!\R.aluOp.ALUOpSRL~q\ & ((!\ShiftLeft0~31_combout\) # (!\R.aluOp.ALUOpSLL~q\))) ) ) ) # ( \R.aluOp.ALUOpSRA~q\ & ( !\ShiftRight0~5_combout\ & ( (!\ShiftRight1~33_combout\ & ((!\ShiftLeft0~31_combout\) # (!\R.aluOp.ALUOpSLL~q\))) ) ) ) # ( 
-- !\R.aluOp.ALUOpSRA~q\ & ( !\ShiftRight0~5_combout\ & ( (!\ShiftLeft0~31_combout\) # (!\R.aluOp.ALUOpSLL~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111001100111100001100000010101010100010001010000010000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpSRL~q\,
	datab => \ALT_INV_ShiftLeft0~31_combout\,
	datac => \ALT_INV_ShiftRight1~33_combout\,
	datad => \ALT_INV_R.aluOp.ALUOpSLL~q\,
	datae => \ALT_INV_R.aluOp.ALUOpSRA~q\,
	dataf => \ALT_INV_ShiftRight0~5_combout\,
	combout => \Selector13~0_combout\);

-- Location: LABCELL_X83_Y4_N27
\Selector13~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector13~2_combout\ = ( !\Selector13~0_combout\ & ( !\R.aluData2\(4) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111000011110000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluData2\(4),
	dataf => \ALT_INV_Selector13~0_combout\,
	combout => \Selector13~2_combout\);

-- Location: LABCELL_X80_Y4_N54
\Comb:vJumpAdr[19]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[19]~0_combout\ = ( \Selector13~1_combout\ & ( \Add3~77_sumout\ & ( (!\Equal4~2_combout\) # ((!\R.aluCalc~q\ & ((\R.aluRes\(19)))) # (\R.aluCalc~q\ & (\Selector13~2_combout\))) ) ) ) # ( !\Selector13~1_combout\ & ( \Add3~77_sumout\ & ( 
-- ((!\Equal4~2_combout\) # (\R.aluCalc~q\)) # (\R.aluRes\(19)) ) ) ) # ( \Selector13~1_combout\ & ( !\Add3~77_sumout\ & ( (\Equal4~2_combout\ & ((!\R.aluCalc~q\ & ((\R.aluRes\(19)))) # (\R.aluCalc~q\ & (\Selector13~2_combout\)))) ) ) ) # ( 
-- !\Selector13~1_combout\ & ( !\Add3~77_sumout\ & ( (\Equal4~2_combout\ & ((\R.aluCalc~q\) # (\R.aluRes\(19)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000111111000000000011010111111111001111111111111100110101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector13~2_combout\,
	datab => \ALT_INV_R.aluRes\(19),
	datac => \ALT_INV_R.aluCalc~q\,
	datad => \ALT_INV_Equal4~2_combout\,
	datae => \ALT_INV_Selector13~1_combout\,
	dataf => \ALT_INV_Add3~77_sumout\,
	combout => \Comb:vJumpAdr[19]~0_combout\);

-- Location: FF_X80_Y4_N55
\R.curPC[19]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[19]~0_combout\,
	asdata => \Add0~69_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(19));

-- Location: LABCELL_X81_Y6_N57
\Add0~77\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~77_sumout\ = SUM(( \R.curPC[21]~DUPLICATE_q\ ) + ( GND ) + ( \Add0~74\ ))
-- \Add0~78\ = CARRY(( \R.curPC[21]~DUPLICATE_q\ ) + ( GND ) + ( \Add0~74\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.curPC[21]~DUPLICATE_q\,
	cin => \Add0~74\,
	sumout => \Add0~77_sumout\,
	cout => \Add0~78\);

-- Location: LABCELL_X81_Y5_N30
\Add0~81\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~81_sumout\ = SUM(( \R.curPC\(22) ) + ( GND ) + ( \Add0~78\ ))
-- \Add0~82\ = CARRY(( \R.curPC\(22) ) + ( GND ) + ( \Add0~78\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.curPC\(22),
	cin => \Add0~78\,
	sumout => \Add0~81_sumout\,
	cout => \Add0~82\);

-- Location: LABCELL_X81_Y5_N33
\Add0~85\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~85_sumout\ = SUM(( \R.curPC\(23) ) + ( GND ) + ( \Add0~82\ ))
-- \Add0~86\ = CARRY(( \R.curPC\(23) ) + ( GND ) + ( \Add0~82\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curPC\(23),
	cin => \Add0~82\,
	sumout => \Add0~85_sumout\,
	cout => \Add0~86\);

-- Location: LABCELL_X81_Y8_N48
\ShiftLeft0~41\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~41_combout\ = ( \R.aluData2\(3) & ( \ShiftLeft0~32_OTERM297\ & ( (!\R.aluData2\(2) & (\ShiftLeft0~24_OTERM293\)) # (\R.aluData2\(2) & ((\ShiftLeft0~16_OTERM287\))) ) ) ) # ( !\R.aluData2\(3) & ( \ShiftLeft0~32_OTERM297\ & ( 
-- (\ShiftLeft0~40_OTERM755\) # (\R.aluData2\(2)) ) ) ) # ( \R.aluData2\(3) & ( !\ShiftLeft0~32_OTERM297\ & ( (!\R.aluData2\(2) & (\ShiftLeft0~24_OTERM293\)) # (\R.aluData2\(2) & ((\ShiftLeft0~16_OTERM287\))) ) ) ) # ( !\R.aluData2\(3) & ( 
-- !\ShiftLeft0~32_OTERM297\ & ( (!\R.aluData2\(2) & \ShiftLeft0~40_OTERM755\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011110000010100110101001100001111111111110101001101010011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~24_OTERM293\,
	datab => \ALT_INV_ShiftLeft0~16_OTERM287\,
	datac => \ALT_INV_R.aluData2\(2),
	datad => \ALT_INV_ShiftLeft0~40_OTERM755\,
	datae => \ALT_INV_R.aluData2\(3),
	dataf => \ALT_INV_ShiftLeft0~32_OTERM297\,
	combout => \ShiftLeft0~41_combout\);

-- Location: LABCELL_X77_Y8_N27
\Selector8~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector8~0_combout\ = ( \R.aluData1\(31) & ( (\R.aluData2\(3) & \R.aluOp.ALUOpSRA~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000011110000000000001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluData2\(3),
	datad => \ALT_INV_R.aluOp.ALUOpSRA~q\,
	dataf => \ALT_INV_R.aluData1\(31),
	combout => \Selector8~0_combout\);

-- Location: LABCELL_X81_Y8_N30
\Selector8~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector8~1_combout\ = ( !\R.aluData2\(4) & ( \R.aluOp.ALUOpSLL~q\ & ( (((\Selector31~0_OTERM349\ & \ShiftRight0~10_combout\)) # (\Selector8~0_combout\)) # (\ShiftLeft0~41_combout\) ) ) ) # ( !\R.aluData2\(4) & ( !\R.aluOp.ALUOpSLL~q\ & ( 
-- ((\Selector31~0_OTERM349\ & \ShiftRight0~10_combout\)) # (\Selector8~0_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100111111000000000000000001011111011111110000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~41_combout\,
	datab => \ALT_INV_Selector31~0_OTERM349\,
	datac => \ALT_INV_Selector8~0_combout\,
	datad => \ALT_INV_ShiftRight0~10_combout\,
	datae => \ALT_INV_R.aluData2\(4),
	dataf => \ALT_INV_R.aluOp.ALUOpSLL~q\,
	combout => \Selector8~1_combout\);

-- Location: MLABCELL_X82_Y4_N6
\Selector8~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector8~2_combout\ = ( \R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( \R.aluOp.ALUOpOr~q\ & ( (!\R.aluData1\(24) & !\R.aluData2\(24)) ) ) ) # ( !\R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( \R.aluOp.ALUOpOr~q\ & ( (!\R.aluData1\(24) & !\R.aluData2\(24)) ) ) ) # ( 
-- \R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( !\R.aluOp.ALUOpOr~q\ & ( (!\R.aluOp.ALUOpXor~DUPLICATE_q\ & ((!\R.aluData1\(24)) # (!\R.aluData2\(24)))) # (\R.aluOp.ALUOpXor~DUPLICATE_q\ & (!\R.aluData1\(24) & !\R.aluData2\(24))) ) ) ) # ( 
-- !\R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( !\R.aluOp.ALUOpOr~q\ & ( (!\R.aluOp.ALUOpXor~DUPLICATE_q\) # (!\R.aluData1\(24) $ (\R.aluData2\(24))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111101010101111111110101010000011110000000000001111000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpXor~DUPLICATE_q\,
	datac => \ALT_INV_R.aluData1\(24),
	datad => \ALT_INV_R.aluData2\(24),
	datae => \ALT_INV_R.aluOp.ALUOpAnd~DUPLICATE_q\,
	dataf => \ALT_INV_R.aluOp.ALUOpOr~q\,
	combout => \Selector8~2_combout\);

-- Location: LABCELL_X81_Y4_N3
\Selector8~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector8~3_combout\ = ( \ShiftLeft0~11_combout\ & ( !\Selector17~0_OTERM391\ & ( (!\Selector12~2_OTERM395\ & \Selector8~2_combout\) ) ) ) # ( !\ShiftLeft0~11_combout\ & ( !\Selector17~0_OTERM391\ & ( \Selector8~2_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111000000001010101000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector12~2_OTERM395\,
	datad => \ALT_INV_Selector8~2_combout\,
	datae => \ALT_INV_ShiftLeft0~11_combout\,
	dataf => \ALT_INV_Selector17~0_OTERM391\,
	combout => \Selector8~3_combout\);

-- Location: LABCELL_X80_Y4_N42
\Comb:vRegWriteData[24]~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[24]~4_combout\ = ( \Selector8~3_combout\ & ( (!\R.aluCalc~q\ & (!\R.aluRes\(24) & (!\R.memToReg~q\))) # (\R.aluCalc~q\ & (((!\Selector8~1_combout\)))) ) ) # ( !\Selector8~3_combout\ & ( (!\R.aluRes\(24) & (!\R.aluCalc~q\ & 
-- !\R.memToReg~q\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000000010000000100000001000000010110011100000001011001110000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluRes\(24),
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_R.memToReg~q\,
	datad => \ALT_INV_Selector8~1_combout\,
	dataf => \ALT_INV_Selector8~3_combout\,
	combout => \Comb:vRegWriteData[24]~4_combout\);

-- Location: LABCELL_X81_Y5_N18
\Comb:vRegWriteData[24]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[24]~2_combout\ = ( \Add1~97_sumout\ & ( \R.curInst\(12) & ( (!\R.memToReg~q\ & (((\R.aluOp.ALUOpAdd~q\)))) # (\R.memToReg~q\ & (!\R.curInst\(14) & (\avm_d_readdata[23]~input_o\))) ) ) ) # ( !\Add1~97_sumout\ & ( \R.curInst\(12) & ( 
-- (!\R.curInst\(14) & (\avm_d_readdata[23]~input_o\ & \R.memToReg~q\)) ) ) ) # ( \Add1~97_sumout\ & ( !\R.curInst\(12) & ( (!\R.memToReg~q\ & ((\R.aluOp.ALUOpAdd~q\))) # (\R.memToReg~q\ & (!\R.curInst\(14))) ) ) ) # ( !\Add1~97_sumout\ & ( !\R.curInst\(12) 
-- & ( (!\R.curInst\(14) & \R.memToReg~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000010101010000011111010101000000000001000100000111100100010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(14),
	datab => \ALT_INV_avm_d_readdata[23]~input_o\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_R.memToReg~q\,
	datae => \ALT_INV_Add1~97_sumout\,
	dataf => \ALT_INV_R.curInst\(12),
	combout => \Comb:vRegWriteData[24]~2_combout\);

-- Location: IOIBUF_X72_Y0_N35
\avm_d_readdata[0]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(0),
	o => \avm_d_readdata[0]~input_o\);

-- Location: LABCELL_X79_Y1_N6
\Comb:vRegWriteData[24]~3_RESYN1104\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[24]~3_RESYN1104_BDD1105\ = ( \avm_d_readdata[0]~input_o\ & ( (!\avm_d_readdata[31]~input_o\ & !\R.curInst\(13)) ) ) # ( !\avm_d_readdata[0]~input_o\ & ( (!\avm_d_readdata[31]~input_o\) # (\R.curInst\(13)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1100110011111111110011001111111111001100000000001100110000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_avm_d_readdata[31]~input_o\,
	datad => \ALT_INV_R.curInst\(13),
	dataf => \ALT_INV_avm_d_readdata[0]~input_o\,
	combout => \Comb:vRegWriteData[24]~3_RESYN1104_BDD1105\);

-- Location: LABCELL_X79_Y1_N12
\Comb:vRegWriteData[24]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[24]~3_combout\ = ( \R.curInst\(13) & ( \R.curInst\(12) & ( \R.memToReg~q\ ) ) ) # ( !\R.curInst\(13) & ( \R.curInst\(12) & ( (\R.memToReg~q\ & ((!\avm_d_readdata[23]~input_o\) # (\R.curInst\(14)))) ) ) ) # ( \R.curInst\(13) & ( 
-- !\R.curInst\(12) & ( (\R.memToReg~q\ & ((\Comb:vRegWriteData[24]~3_RESYN1104_BDD1105\) # (\R.curInst\(14)))) ) ) ) # ( !\R.curInst\(13) & ( !\R.curInst\(12) & ( (\R.memToReg~q\ & ((\Comb:vRegWriteData[24]~3_RESYN1104_BDD1105\) # (\R.curInst\(14)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100110011000000110011001100100011001000110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_avm_d_readdata[23]~input_o\,
	datab => \ALT_INV_R.memToReg~q\,
	datac => \ALT_INV_R.curInst\(14),
	datad => \ALT_INV_Comb:vRegWriteData[24]~3_RESYN1104_BDD1105\,
	datae => \ALT_INV_R.curInst\(13),
	dataf => \ALT_INV_R.curInst\(12),
	combout => \Comb:vRegWriteData[24]~3_combout\);

-- Location: LABCELL_X81_Y5_N12
\Comb:vRegWriteData[24]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[24]~0_combout\ = ( !\Comb:vRegWriteData[24]~3_combout\ & ( \Add2~97_sumout\ & ( (!\Comb:vRegWriteData[24]~4_combout\) # ((\R.aluCalc~q\ & ((\Comb:vRegWriteData[24]~2_combout\) # (\R.aluOp.ALUOpSub~q\)))) ) ) ) # ( 
-- !\Comb:vRegWriteData[24]~3_combout\ & ( !\Add2~97_sumout\ & ( (!\Comb:vRegWriteData[24]~4_combout\) # ((\Comb:vRegWriteData[24]~2_combout\ & \R.aluCalc~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010101010101111000000000000000010101010101111110000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Comb:vRegWriteData[24]~4_combout\,
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_Comb:vRegWriteData[24]~2_combout\,
	datad => \ALT_INV_R.aluCalc~q\,
	datae => \ALT_INV_Comb:vRegWriteData[24]~3_combout\,
	dataf => \ALT_INV_Add2~97_sumout\,
	combout => \Comb:vRegWriteData[24]~0_combout\);

-- Location: FF_X81_Y5_N38
\R.regWriteData[24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Add0~89_sumout\,
	asdata => \Comb:vRegWriteData[24]~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(24));

-- Location: FF_X68_Y1_N38
\RegFile[29][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(24),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][24]~q\);

-- Location: FF_X67_Y1_N56
\RegFile[31][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(24),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][24]~q\);

-- Location: LABCELL_X66_Y3_N45
\RegFile[30][24]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[30][24]~feeder_combout\ = ( \R.regWriteData\(24) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(24),
	combout => \RegFile[30][24]~feeder_combout\);

-- Location: FF_X66_Y3_N46
\RegFile[30][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[30][24]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][24]~q\);

-- Location: LABCELL_X67_Y1_N30
\RegFile[25][24]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[25][24]~feeder_combout\ = ( \R.regWriteData\(24) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(24),
	combout => \RegFile[25][24]~feeder_combout\);

-- Location: FF_X67_Y1_N32
\RegFile[25][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[25][24]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][24]~q\);

-- Location: FF_X67_Y1_N44
\RegFile[27][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(24),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][24]~q\);

-- Location: FF_X67_Y2_N52
\RegFile[26][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(24),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][24]~q\);

-- Location: MLABCELL_X59_Y2_N0
\RegFile[24][24]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[24][24]~feeder_combout\ = ( \R.regWriteData\(24) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(24),
	combout => \RegFile[24][24]~feeder_combout\);

-- Location: FF_X59_Y2_N1
\RegFile[24][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[24][24]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][24]~q\);

-- Location: LABCELL_X68_Y1_N12
\Mux98~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux98~22_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[24][24]~q\))) # (\R.curInst\(20) & (\RegFile[25][24]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[26][24]~q\))) # (\R.curInst\(20) & (\RegFile[27][24]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[25][24]~q\,
	datab => \ALT_INV_RegFile[27][24]~q\,
	datac => \ALT_INV_RegFile[26][24]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][24]~q\,
	combout => \Mux98~22_combout\);

-- Location: FF_X66_Y3_N4
\RegFile[28][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(24),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][24]~q\);

-- Location: LABCELL_X68_Y1_N36
\Mux98~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux98~9_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux98~22_combout\)))) # (\R.curInst\(22) & ((!\Mux98~22_combout\ & ((\RegFile[28][24]~q\))) # (\Mux98~22_combout\ & (\RegFile[29][24]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux98~22_combout\)))) # (\R.curInst\(22) & ((!\Mux98~22_combout\ & ((\RegFile[30][24]~q\))) # (\Mux98~22_combout\ & (\RegFile[31][24]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[29][24]~q\,
	datab => \ALT_INV_RegFile[31][24]~q\,
	datac => \ALT_INV_RegFile[30][24]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux98~22_combout\,
	datag => \ALT_INV_RegFile[28][24]~q\,
	combout => \Mux98~9_combout\);

-- Location: FF_X67_Y3_N20
\RegFile[3][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(24),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][24]~q\);

-- Location: LABCELL_X60_Y5_N12
\RegFile[2][24]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[2][24]~feeder_combout\ = ( \R.regWriteData\(24) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(24),
	combout => \RegFile[2][24]~feeder_combout\);

-- Location: FF_X60_Y5_N13
\RegFile[2][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[2][24]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][24]~q\);

-- Location: LABCELL_X60_Y3_N30
\RegFile[5][24]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[5][24]~feeder_combout\ = ( \R.regWriteData\(24) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(24),
	combout => \RegFile[5][24]~feeder_combout\);

-- Location: FF_X60_Y3_N31
\RegFile[5][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[5][24]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][24]~q\);

-- Location: FF_X67_Y3_N49
\RegFile[7][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(24),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][24]~q\);

-- Location: FF_X67_Y3_N8
\RegFile[6][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(24),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][24]~q\);

-- Location: LABCELL_X60_Y3_N24
\RegFile[4][24]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[4][24]~feeder_combout\ = ( \R.regWriteData\(24) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(24),
	combout => \RegFile[4][24]~feeder_combout\);

-- Location: FF_X60_Y3_N25
\RegFile[4][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[4][24]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][24]~q\);

-- Location: LABCELL_X62_Y3_N6
\Mux98~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux98~0_combout\ = ( \R.curInst\(21) & ( \R.curInst\(20) & ( \RegFile[7][24]~q\ ) ) ) # ( !\R.curInst\(21) & ( \R.curInst\(20) & ( \RegFile[5][24]~q\ ) ) ) # ( \R.curInst\(21) & ( !\R.curInst\(20) & ( \RegFile[6][24]~q\ ) ) ) # ( !\R.curInst\(21) & ( 
-- !\R.curInst\(20) & ( \RegFile[4][24]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111000011110000111101010101010101010011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[5][24]~q\,
	datab => \ALT_INV_RegFile[7][24]~q\,
	datac => \ALT_INV_RegFile[6][24]~q\,
	datad => \ALT_INV_RegFile[4][24]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	combout => \Mux98~0_combout\);

-- Location: FF_X61_Y5_N49
\RegFile[1][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(24),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][24]~q\);

-- Location: LABCELL_X60_Y5_N48
\Mux98~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux98~26_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (\R.curInst\(20) & (\RegFile[1][24]~q\))) # (\R.curInst\(22) & (((\Mux98~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (((\RegFile[2][24]~q\)))) # 
-- (\R.curInst\(20) & (\RegFile[3][24]~q\)))) # (\R.curInst\(22) & ((((\Mux98~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000000000111010000000000000011111111110001110111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][24]~q\,
	datab => \ALT_INV_R.curInst\(20),
	datac => \ALT_INV_RegFile[2][24]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux98~0_combout\,
	datag => \ALT_INV_RegFile[1][24]~q\,
	combout => \Mux98~26_combout\);

-- Location: FF_X62_Y2_N56
\RegFile[13][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(24),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][24]~q\);

-- Location: FF_X70_Y1_N32
\RegFile[15][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(24),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][24]~q\);

-- Location: FF_X65_Y5_N28
\RegFile[14][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(24),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][24]~q\);

-- Location: FF_X70_Y2_N49
\RegFile[9][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(24),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][24]~q\);

-- Location: FF_X64_Y3_N19
\RegFile[10][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(24),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][24]~q\);

-- Location: FF_X70_Y1_N26
\RegFile[11][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(24),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][24]~q\);

-- Location: LABCELL_X66_Y5_N21
\RegFile[8][24]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[8][24]~feeder_combout\ = ( \R.regWriteData\(24) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(24),
	combout => \RegFile[8][24]~feeder_combout\);

-- Location: FF_X66_Y5_N22
\RegFile[8][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[8][24]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][24]~q\);

-- Location: LABCELL_X66_Y2_N54
\Mux98~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux98~14_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[8][24]~q\))) # (\R.curInst\(20) & (\RegFile[9][24]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & (\RegFile[10][24]~q\)) # (\R.curInst\(20) & ((\RegFile[11][24]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][24]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[10][24]~q\,
	datad => \ALT_INV_RegFile[11][24]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][24]~q\,
	combout => \Mux98~14_combout\);

-- Location: LABCELL_X62_Y2_N6
\RegFile[12][24]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[12][24]~feeder_combout\ = ( \R.regWriteData\(24) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(24),
	combout => \RegFile[12][24]~feeder_combout\);

-- Location: FF_X62_Y2_N8
\RegFile[12][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[12][24]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][24]~q\);

-- Location: LABCELL_X62_Y5_N0
\Mux98~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux98~1_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux98~14_combout\)))) # (\R.curInst\(22) & ((!\Mux98~14_combout\ & ((\RegFile[12][24]~q\))) # (\Mux98~14_combout\ & (\RegFile[13][24]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux98~14_combout\)))) # (\R.curInst\(22) & ((!\Mux98~14_combout\ & ((\RegFile[14][24]~q\))) # (\Mux98~14_combout\ & (\RegFile[15][24]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][24]~q\,
	datab => \ALT_INV_RegFile[15][24]~q\,
	datac => \ALT_INV_RegFile[14][24]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux98~14_combout\,
	datag => \ALT_INV_RegFile[12][24]~q\,
	combout => \Mux98~1_combout\);

-- Location: FF_X70_Y1_N2
\RegFile[23][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(24),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][24]~q\);

-- Location: FF_X61_Y6_N22
\RegFile[21][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(24),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][24]~q\);

-- Location: FF_X61_Y6_N49
\RegFile[22][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(24),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][24]~q\);

-- Location: FF_X64_Y2_N20
\RegFile[17][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(24),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][24]~q\);

-- Location: LABCELL_X64_Y2_N54
\RegFile[19][24]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[19][24]~feeder_combout\ = ( \R.regWriteData\(24) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(24),
	combout => \RegFile[19][24]~feeder_combout\);

-- Location: FF_X64_Y2_N55
\RegFile[19][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[19][24]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][24]~q\);

-- Location: MLABCELL_X59_Y3_N3
\RegFile[18][24]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[18][24]~feeder_combout\ = ( \R.regWriteData\(24) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(24),
	combout => \RegFile[18][24]~feeder_combout\);

-- Location: FF_X59_Y3_N4
\RegFile[18][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][24]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][24]~q\);

-- Location: FF_X64_Y1_N35
\RegFile[16][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(24),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][24]~q\);

-- Location: LABCELL_X64_Y2_N18
\Mux98~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux98~18_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[16][24]~q\))) # (\R.curInst\(20) & (\RegFile[17][24]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[18][24]~q\))) # (\R.curInst\(20) & (\RegFile[19][24]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[17][24]~q\,
	datab => \ALT_INV_RegFile[19][24]~q\,
	datac => \ALT_INV_RegFile[18][24]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][24]~q\,
	combout => \Mux98~18_combout\);

-- Location: MLABCELL_X59_Y3_N27
\RegFile[20][24]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[20][24]~feeder_combout\ = ( \R.regWriteData\(24) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(24),
	combout => \RegFile[20][24]~feeder_combout\);

-- Location: FF_X59_Y3_N28
\RegFile[20][24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[20][24]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][24]~q\);

-- Location: LABCELL_X61_Y3_N24
\Mux98~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux98~5_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux98~18_combout\)))) # (\R.curInst\(22) & ((!\Mux98~18_combout\ & ((\RegFile[20][24]~q\))) # (\Mux98~18_combout\ & (\RegFile[21][24]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux98~18_combout\)))) # (\R.curInst\(22) & ((!\Mux98~18_combout\ & ((\RegFile[22][24]~q\))) # (\Mux98~18_combout\ & (\RegFile[23][24]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[23][24]~q\,
	datab => \ALT_INV_RegFile[21][24]~q\,
	datac => \ALT_INV_RegFile[22][24]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux98~18_combout\,
	datag => \ALT_INV_RegFile[20][24]~q\,
	combout => \Mux98~5_combout\);

-- Location: LABCELL_X61_Y5_N45
\Mux98~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux98~13_combout\ = ( \Mux98~1_combout\ & ( \Mux98~5_combout\ & ( (!\R.curInst\(24) & (((\R.curInst\(23)) # (\Mux98~26_combout\)))) # (\R.curInst\(24) & (((!\R.curInst\(23))) # (\Mux98~9_combout\))) ) ) ) # ( !\Mux98~1_combout\ & ( \Mux98~5_combout\ & ( 
-- (!\R.curInst\(24) & (((\Mux98~26_combout\ & !\R.curInst\(23))))) # (\R.curInst\(24) & (((!\R.curInst\(23))) # (\Mux98~9_combout\))) ) ) ) # ( \Mux98~1_combout\ & ( !\Mux98~5_combout\ & ( (!\R.curInst\(24) & (((\R.curInst\(23)) # (\Mux98~26_combout\)))) # 
-- (\R.curInst\(24) & (\Mux98~9_combout\ & ((\R.curInst\(23))))) ) ) ) # ( !\Mux98~1_combout\ & ( !\Mux98~5_combout\ & ( (!\R.curInst\(24) & (((\Mux98~26_combout\ & !\R.curInst\(23))))) # (\R.curInst\(24) & (\Mux98~9_combout\ & ((\R.curInst\(23))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101000010001000010101011101101011111000100010101111110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(24),
	datab => \ALT_INV_Mux98~9_combout\,
	datac => \ALT_INV_Mux98~26_combout\,
	datad => \ALT_INV_R.curInst\(23),
	datae => \ALT_INV_Mux98~1_combout\,
	dataf => \ALT_INV_Mux98~5_combout\,
	combout => \Mux98~13_combout\);

-- Location: LABCELL_X75_Y5_N3
\NxR.aluData2[24]~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[24]~26_combout\ = ( \Equal4~1_combout\ & ( \Mux98~13_combout\ & ( (!\vAluSrc2~1_combout\) # (\Mux130~0_combout\) ) ) ) # ( !\Equal4~1_combout\ & ( \Mux98~13_combout\ & ( !\vAluSrc2~1_combout\ ) ) ) # ( \Equal4~1_combout\ & ( 
-- !\Mux98~13_combout\ & ( (\Mux130~0_combout\ & \vAluSrc2~1_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000100010001000111001100110011001101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux130~0_combout\,
	datab => \ALT_INV_vAluSrc2~1_combout\,
	datae => \ALT_INV_Equal4~1_combout\,
	dataf => \ALT_INV_Mux98~13_combout\,
	combout => \NxR.aluData2[24]~26_combout\);

-- Location: FF_X75_Y5_N4
\R.aluData2[24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR.aluData2[24]~26_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData2\(24));

-- Location: LABCELL_X80_Y4_N36
\Selector8~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector8~4_combout\ = ( \Add1~97_sumout\ & ( \Selector8~3_combout\ & ( (((\R.aluOp.ALUOpSub~q\ & \Add2~97_sumout\)) # (\Selector8~1_combout\)) # (\R.aluOp.ALUOpAdd~q\) ) ) ) # ( !\Add1~97_sumout\ & ( \Selector8~3_combout\ & ( ((\R.aluOp.ALUOpSub~q\ & 
-- \Add2~97_sumout\)) # (\Selector8~1_combout\) ) ) ) # ( \Add1~97_sumout\ & ( !\Selector8~3_combout\ ) ) # ( !\Add1~97_sumout\ & ( !\Selector8~3_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111111111111111111100000101111111110011011111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datab => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datac => \ALT_INV_Add2~97_sumout\,
	datad => \ALT_INV_Selector8~1_combout\,
	datae => \ALT_INV_Add1~97_sumout\,
	dataf => \ALT_INV_Selector8~3_combout\,
	combout => \Selector8~4_combout\);

-- Location: LABCELL_X80_Y4_N18
\Comb:vJumpAdr[24]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[24]~0_combout\ = ( \Add3~97_sumout\ & ( (!\Equal4~2_combout\) # ((!\R.aluCalc~q\ & ((\R.aluRes\(24)))) # (\R.aluCalc~q\ & (\Selector8~4_combout\))) ) ) # ( !\Add3~97_sumout\ & ( (\Equal4~2_combout\ & ((!\R.aluCalc~q\ & ((\R.aluRes\(24)))) # 
-- (\R.aluCalc~q\ & (\Selector8~4_combout\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000011101000000000001110111111111000111011111111100011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector8~4_combout\,
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_R.aluRes\(24),
	datad => \ALT_INV_Equal4~2_combout\,
	dataf => \ALT_INV_Add3~97_sumout\,
	combout => \Comb:vJumpAdr[24]~0_combout\);

-- Location: FF_X80_Y4_N19
\R.curPC[24]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[24]~0_combout\,
	asdata => \Add0~89_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(24));

-- Location: LABCELL_X70_Y1_N24
\Mux66~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux66~14_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[8][24]~q\))) # (\R.curInst\(15) & (\RegFile[9][24]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[10][24]~q\))) # (\R.curInst\(15) & (\RegFile[11][24]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[11][24]~q\,
	datab => \ALT_INV_RegFile[9][24]~q\,
	datac => \ALT_INV_RegFile[10][24]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][24]~q\,
	combout => \Mux66~14_combout\);

-- Location: LABCELL_X70_Y1_N30
\Mux66~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux66~1_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux66~14_combout\))))) # (\R.curInst\(17) & (((!\Mux66~14_combout\ & ((\RegFile[12][24]~q\))) # (\Mux66~14_combout\ & (\RegFile[13][24]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux66~14_combout\)))) # (\R.curInst\(17) & ((!\Mux66~14_combout\ & (\RegFile[14][24]~q\)) # (\Mux66~14_combout\ & ((\RegFile[15][24]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][24]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[14][24]~q\,
	datad => \ALT_INV_RegFile[15][24]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux66~14_combout\,
	datag => \ALT_INV_RegFile[12][24]~q\,
	combout => \Mux66~1_combout\);

-- Location: LABCELL_X67_Y1_N42
\Mux66~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux66~22_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & (\RegFile[24][24]~q\)) # (\R.curInst\(15) & ((\RegFile[25][24]~q\)))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & ((\RegFile[26][24]~q\))) # (\R.curInst\(15) & (\RegFile[27][24]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001010101111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[27][24]~q\,
	datac => \ALT_INV_RegFile[26][24]~q\,
	datad => \ALT_INV_RegFile[25][24]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][24]~q\,
	combout => \Mux66~22_combout\);

-- Location: LABCELL_X67_Y1_N54
\Mux66~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux66~9_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux66~22_combout\)))) # (\R.curInst\(17) & ((!\Mux66~22_combout\ & ((\RegFile[28][24]~q\))) # (\Mux66~22_combout\ & (\RegFile[29][24]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux66~22_combout\)))) # (\R.curInst\(17) & ((!\Mux66~22_combout\ & ((\RegFile[30][24]~q\))) # (\Mux66~22_combout\ & (\RegFile[31][24]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][24]~q\,
	datab => \ALT_INV_RegFile[29][24]~q\,
	datac => \ALT_INV_RegFile[30][24]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux66~22_combout\,
	datag => \ALT_INV_RegFile[28][24]~q\,
	combout => \Mux66~9_combout\);

-- Location: LABCELL_X64_Y2_N30
\Mux66~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux66~18_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[16][24]~q\))) # (\R.curInst\(15) & (\RegFile[17][24]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[18][24]~q\))) # (\R.curInst\(15) & (\RegFile[19][24]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[17][24]~q\,
	datab => \ALT_INV_RegFile[19][24]~q\,
	datac => \ALT_INV_RegFile[18][24]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][24]~q\,
	combout => \Mux66~18_combout\);

-- Location: LABCELL_X70_Y1_N0
\Mux66~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux66~5_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux66~18_combout\))))) # (\R.curInst\(17) & (((!\Mux66~18_combout\ & ((\RegFile[20][24]~q\))) # (\Mux66~18_combout\ & (\RegFile[21][24]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux66~18_combout\)))) # (\R.curInst\(17) & ((!\Mux66~18_combout\ & (\RegFile[22][24]~q\)) # (\Mux66~18_combout\ & ((\RegFile[23][24]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][24]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[22][24]~q\,
	datad => \ALT_INV_RegFile[23][24]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux66~18_combout\,
	datag => \ALT_INV_RegFile[20][24]~q\,
	combout => \Mux66~5_combout\);

-- Location: LABCELL_X67_Y3_N48
\Mux66~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux66~0_combout\ = ( \RegFile[7][24]~q\ & ( \R.curInst\(15) & ( (\RegFile[5][24]~q\) # (\R.curInst\(16)) ) ) ) # ( !\RegFile[7][24]~q\ & ( \R.curInst\(15) & ( (!\R.curInst\(16) & \RegFile[5][24]~q\) ) ) ) # ( \RegFile[7][24]~q\ & ( !\R.curInst\(15) & ( 
-- (!\R.curInst\(16) & ((\RegFile[4][24]~q\))) # (\R.curInst\(16) & (\RegFile[6][24]~q\)) ) ) ) # ( !\RegFile[7][24]~q\ & ( !\R.curInst\(15) & ( (!\R.curInst\(16) & ((\RegFile[4][24]~q\))) # (\R.curInst\(16) & (\RegFile[6][24]~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001101100011011000110110001101100000000101010100101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(16),
	datab => \ALT_INV_RegFile[6][24]~q\,
	datac => \ALT_INV_RegFile[4][24]~q\,
	datad => \ALT_INV_RegFile[5][24]~q\,
	datae => \ALT_INV_RegFile[7][24]~q\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux66~0_combout\);

-- Location: LABCELL_X67_Y3_N30
\Mux66~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux66~26_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (\RegFile[1][24]~q\ & (\R.curInst\(15)))) # (\R.curInst\(17) & (((\Mux66~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & ((!\R.curInst\(15) & (((\RegFile[2][24]~q\)))) # 
-- (\R.curInst\(15) & (\RegFile[3][24]~q\)))) # (\R.curInst\(17) & ((((\Mux66~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001100000011000100010000110011001111110011111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][24]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[2][24]~q\,
	datad => \ALT_INV_R.curInst\(15),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux66~0_combout\,
	datag => \ALT_INV_RegFile[1][24]~q\,
	combout => \Mux66~26_combout\);

-- Location: LABCELL_X70_Y1_N48
\Mux66~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux66~13_combout\ = ( \Mux66~5_combout\ & ( \Mux66~26_combout\ & ( (!\R.curInst\(18)) # ((!\R.curInst\(19) & (\Mux66~1_combout\)) # (\R.curInst\(19) & ((\Mux66~9_combout\)))) ) ) ) # ( !\Mux66~5_combout\ & ( \Mux66~26_combout\ & ( (!\R.curInst\(19) & 
-- ((!\R.curInst\(18)) # ((\Mux66~1_combout\)))) # (\R.curInst\(19) & (\R.curInst\(18) & ((\Mux66~9_combout\)))) ) ) ) # ( \Mux66~5_combout\ & ( !\Mux66~26_combout\ & ( (!\R.curInst\(19) & (\R.curInst\(18) & (\Mux66~1_combout\))) # (\R.curInst\(19) & 
-- ((!\R.curInst\(18)) # ((\Mux66~9_combout\)))) ) ) ) # ( !\Mux66~5_combout\ & ( !\Mux66~26_combout\ & ( (\R.curInst\(18) & ((!\R.curInst\(19) & (\Mux66~1_combout\)) # (\R.curInst\(19) & ((\Mux66~9_combout\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001000010011010001100101011110001010100110111100111011011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(19),
	datab => \ALT_INV_R.curInst\(18),
	datac => \ALT_INV_Mux66~1_combout\,
	datad => \ALT_INV_Mux66~9_combout\,
	datae => \ALT_INV_Mux66~5_combout\,
	dataf => \ALT_INV_Mux66~26_combout\,
	combout => \Mux66~13_combout\);

-- Location: LABCELL_X74_Y3_N21
\Mux230~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux230~0_combout\ = ( \Mux66~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC\(24)))) ) ) # ( !\Mux66~13_combout\ & ( (\R.curPC\(24) & (\vAluSrc1~2_combout\ & !\vAluSrc1~1_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100000000000100010000000011011101000000001101110100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curPC\(24),
	datab => \ALT_INV_vAluSrc1~2_combout\,
	datad => \ALT_INV_vAluSrc1~1_combout\,
	dataf => \ALT_INV_Mux66~13_combout\,
	combout => \Mux230~0_combout\);

-- Location: LABCELL_X74_Y3_N3
\ShiftRight1~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~26_combout\ = ( \NxR.aluData2[0]~16_combout\ & ( \Mux229~0_combout\ & ( (\NxR.aluData2[1]~17_combout\) # (\Mux231~0_combout\) ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( \Mux229~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & 
-- ((\Mux232~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux230~0_combout\)) ) ) ) # ( \NxR.aluData2[0]~16_combout\ & ( !\Mux229~0_combout\ & ( (\Mux231~0_combout\ & !\NxR.aluData2[1]~17_combout\) ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( 
-- !\Mux229~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((\Mux232~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux230~0_combout\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010111110101001100000011000000000101111101010011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux230~0_combout\,
	datab => \ALT_INV_Mux231~0_combout\,
	datac => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datad => \ALT_INV_Mux232~0_combout\,
	datae => \ALT_INV_NxR.aluData2[0]~16_combout\,
	dataf => \ALT_INV_Mux229~0_combout\,
	combout => \ShiftRight1~26_combout\);

-- Location: FF_X74_Y3_N4
\ShiftRight1~26_NEW_REG36\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~26_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~26_OTERM37\);

-- Location: LABCELL_X73_Y6_N57
\ShiftRight1~28\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~28_combout\ = ( \Mux224~0_combout\ & ( ((!\NxR.aluData2[0]~16_combout\ & !\NxR.aluData2[1]~17_combout\)) # (\Mux223~0_combout\) ) ) # ( !\Mux224~0_combout\ & ( (\Mux223~0_combout\ & ((\NxR.aluData2[1]~17_combout\) # 
-- (\NxR.aluData2[0]~16_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100001111000001010000111110101111000011111010111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datac => \ALT_INV_Mux223~0_combout\,
	datad => \ALT_INV_NxR.aluData2[1]~17_combout\,
	dataf => \ALT_INV_Mux224~0_combout\,
	combout => \ShiftRight1~28_combout\);

-- Location: FF_X73_Y6_N58
\ShiftRight1~28_NEW_REG22\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~28_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~28_OTERM23\);

-- Location: MLABCELL_X82_Y6_N42
\ShiftRight1~43\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~43_combout\ = ( \R.aluData2\(2) & ( \R.aluData1\(31) & ( (\ShiftRight1~27_OTERM19\) # (\R.aluData2\(3)) ) ) ) # ( !\R.aluData2\(2) & ( \R.aluData1\(31) & ( (!\R.aluData2\(3) & (\ShiftRight1~26_OTERM37\)) # (\R.aluData2\(3) & 
-- ((\ShiftRight1~28_OTERM23\))) ) ) ) # ( \R.aluData2\(2) & ( !\R.aluData1\(31) & ( (!\R.aluData2\(3) & \ShiftRight1~27_OTERM19\) ) ) ) # ( !\R.aluData2\(2) & ( !\R.aluData1\(31) & ( (!\R.aluData2\(3) & (\ShiftRight1~26_OTERM37\)) # (\R.aluData2\(3) & 
-- ((\ShiftRight1~28_OTERM23\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100011101000111000000001100110001000111010001110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~26_OTERM37\,
	datab => \ALT_INV_R.aluData2\(3),
	datac => \ALT_INV_ShiftRight1~28_OTERM23\,
	datad => \ALT_INV_ShiftRight1~27_OTERM19\,
	datae => \ALT_INV_R.aluData2\(2),
	dataf => \ALT_INV_R.aluData1\(31),
	combout => \ShiftRight1~43_combout\);

-- Location: LABCELL_X83_Y6_N9
\Selector26~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector26~4_combout\ = ( \Selector26~0_combout\ ) # ( !\Selector26~0_combout\ & ( (!\Selector26~3_combout\) # ((\Selector31~6_OTERM381\ & \ShiftRight1~43_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111100000101111111110000010111111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector31~6_OTERM381\,
	datac => \ALT_INV_ShiftRight1~43_combout\,
	datad => \ALT_INV_Selector26~3_combout\,
	dataf => \ALT_INV_Selector26~0_combout\,
	combout => \Selector26~4_combout\);

-- Location: FF_X83_Y6_N10
\R.aluRes[6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector26~4_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(6));

-- Location: LABCELL_X80_Y6_N12
\vAluRes~6_RESYN1072\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~6_RESYN1072_BDD1073\ = ( \ShiftRight1~43_combout\ & ( ((\Add2~25_sumout\ & \R.aluOp.ALUOpSub~q\)) # (\Selector31~6_OTERM381\) ) ) # ( !\ShiftRight1~43_combout\ & ( (\Add2~25_sumout\ & \R.aluOp.ALUOpSub~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000001111000000000000111100110011001111110011001100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Selector31~6_OTERM381\,
	datac => \ALT_INV_Add2~25_sumout\,
	datad => \ALT_INV_R.aluOp.ALUOpSub~q\,
	dataf => \ALT_INV_ShiftRight1~43_combout\,
	combout => \vAluRes~6_RESYN1072_BDD1073\);

-- Location: LABCELL_X80_Y6_N30
\vAluRes~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~6_combout\ = ( \Add1~25_sumout\ & ( \Selector26~3_combout\ & ( (!\R.aluCalc~q\ & (((\R.aluRes\(6))))) # (\R.aluCalc~q\ & (((\vAluRes~6_RESYN1072_BDD1073\)) # (\R.aluOp.ALUOpAdd~q\))) ) ) ) # ( !\Add1~25_sumout\ & ( \Selector26~3_combout\ & ( 
-- (!\R.aluCalc~q\ & (\R.aluRes\(6))) # (\R.aluCalc~q\ & ((\vAluRes~6_RESYN1072_BDD1073\))) ) ) ) # ( \Add1~25_sumout\ & ( !\Selector26~3_combout\ & ( (\R.aluCalc~q\) # (\R.aluRes\(6)) ) ) ) # ( !\Add1~25_sumout\ & ( !\Selector26~3_combout\ & ( 
-- (\R.aluCalc~q\) # (\R.aluRes\(6)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011111100111111001111110011111100110000001111110011010100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datab => \ALT_INV_R.aluRes\(6),
	datac => \ALT_INV_R.aluCalc~q\,
	datad => \ALT_INV_vAluRes~6_RESYN1072_BDD1073\,
	datae => \ALT_INV_Add1~25_sumout\,
	dataf => \ALT_INV_Selector26~3_combout\,
	combout => \vAluRes~6_combout\);

-- Location: MLABCELL_X84_Y5_N48
\Comb:vJumpAdr[6]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[6]~0_combout\ = ( \Equal4~2_combout\ & ( \Add3~25_sumout\ & ( \vAluRes~6_combout\ ) ) ) # ( !\Equal4~2_combout\ & ( \Add3~25_sumout\ ) ) # ( \Equal4~2_combout\ & ( !\Add3~25_sumout\ & ( \vAluRes~6_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000111111111111111111110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_vAluRes~6_combout\,
	datae => \ALT_INV_Equal4~2_combout\,
	dataf => \ALT_INV_Add3~25_sumout\,
	combout => \Comb:vJumpAdr[6]~0_combout\);

-- Location: FF_X84_Y5_N49
\R.curPC[6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[6]~0_combout\,
	asdata => \Add0~17_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(6));

-- Location: LABCELL_X67_Y7_N24
\Mux84~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux84~0_combout\ = ( \RegFile[7][6]~q\ & ( \R.curInst\(15) & ( (\RegFile[5][6]~q\) # (\R.curInst\(16)) ) ) ) # ( !\RegFile[7][6]~q\ & ( \R.curInst\(15) & ( (!\R.curInst\(16) & \RegFile[5][6]~q\) ) ) ) # ( \RegFile[7][6]~q\ & ( !\R.curInst\(15) & ( 
-- (!\R.curInst\(16) & (\RegFile[4][6]~q\)) # (\R.curInst\(16) & ((\RegFile[6][6]~q\))) ) ) ) # ( !\RegFile[7][6]~q\ & ( !\R.curInst\(15) & ( (!\R.curInst\(16) & (\RegFile[4][6]~q\)) # (\R.curInst\(16) & ((\RegFile[6][6]~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101001011111000010100101111100100010001000100111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(16),
	datab => \ALT_INV_RegFile[5][6]~q\,
	datac => \ALT_INV_RegFile[4][6]~q\,
	datad => \ALT_INV_RegFile[6][6]~q\,
	datae => \ALT_INV_RegFile[7][6]~q\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux84~0_combout\);

-- Location: LABCELL_X67_Y7_N0
\Mux84~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux84~26_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (\RegFile[1][6]~q\ & (\R.curInst\(15)))) # (\R.curInst\(17) & (((\Mux84~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & ((!\R.curInst\(15) & (((\RegFile[2][6]~q\)))) # 
-- (\R.curInst\(15) & (\RegFile[3][6]~q\)))) # (\R.curInst\(17) & ((((\Mux84~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001100000011000100010000110011001111110011111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][6]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[2][6]~q\,
	datad => \ALT_INV_R.curInst\(15),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux84~0_combout\,
	datag => \ALT_INV_RegFile[1][6]~q\,
	combout => \Mux84~26_combout\);

-- Location: LABCELL_X61_Y7_N0
\Mux84~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux84~22_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[24][6]~q\))) # (\R.curInst\(15) & (\RegFile[25][6]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[26][6]~q\))) # (\R.curInst\(15) & (\RegFile[27][6]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[27][6]~q\,
	datab => \ALT_INV_RegFile[25][6]~q\,
	datac => \ALT_INV_RegFile[26][6]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][6]~q\,
	combout => \Mux84~22_combout\);

-- Location: LABCELL_X62_Y7_N48
\Mux84~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux84~9_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux84~22_combout\)))) # (\R.curInst\(17) & ((!\Mux84~22_combout\ & ((\RegFile[28][6]~q\))) # (\Mux84~22_combout\ & (\RegFile[29][6]~q\))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) 
-- & (((\Mux84~22_combout\)))) # (\R.curInst\(17) & ((!\Mux84~22_combout\ & ((\RegFile[30][6]~q\))) # (\Mux84~22_combout\ & (\RegFile[31][6]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][6]~q\,
	datab => \ALT_INV_RegFile[29][6]~q\,
	datac => \ALT_INV_RegFile[30][6]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux84~22_combout\,
	datag => \ALT_INV_RegFile[28][6]~q\,
	combout => \Mux84~9_combout\);

-- Location: LABCELL_X64_Y7_N12
\Mux84~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux84~18_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & (\RegFile[16][6]~q\)) # (\R.curInst\(15) & ((\RegFile[17][6]~q\))))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & ((\RegFile[18][6]~q\))) # (\R.curInst\(15) & (\RegFile[19][6]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110000110011111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[19][6]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[18][6]~q\,
	datad => \ALT_INV_RegFile[17][6]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][6]~q\,
	combout => \Mux84~18_combout\);

-- Location: LABCELL_X64_Y7_N30
\Mux84~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux84~5_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux84~18_combout\))))) # (\R.curInst\(17) & (((!\Mux84~18_combout\ & ((\RegFile[20][6]~q\))) # (\Mux84~18_combout\ & (\RegFile[21][6]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux84~18_combout\)))) # (\R.curInst\(17) & ((!\Mux84~18_combout\ & (\RegFile[22][6]~q\)) # (\Mux84~18_combout\ & ((\RegFile[23][6]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][6]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[22][6]~q\,
	datad => \ALT_INV_RegFile[23][6]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux84~18_combout\,
	datag => \ALT_INV_RegFile[20][6]~q\,
	combout => \Mux84~5_combout\);

-- Location: FF_X61_Y7_N13
\RegFile[14][6]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(6),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][6]~DUPLICATE_q\);

-- Location: MLABCELL_X65_Y3_N30
\Mux84~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux84~14_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[8][6]~q\))) # (\R.curInst\(15) & (\RegFile[9][6]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & (\RegFile[10][6]~q\)) # (\R.curInst\(15) & ((\RegFile[11][6]~q\)))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001110111011101110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[9][6]~q\,
	datac => \ALT_INV_RegFile[10][6]~q\,
	datad => \ALT_INV_RegFile[11][6]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][6]~q\,
	combout => \Mux84~14_combout\);

-- Location: LABCELL_X66_Y7_N24
\Mux84~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux84~1_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux84~14_combout\)))) # (\R.curInst\(17) & ((!\Mux84~14_combout\ & (\RegFile[12][6]~q\)) # (\Mux84~14_combout\ & ((\RegFile[13][6]~q\)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- ((((\Mux84~14_combout\))))) # (\R.curInst\(17) & (((!\Mux84~14_combout\ & ((\RegFile[14][6]~DUPLICATE_q\))) # (\Mux84~14_combout\ & (\RegFile[15][6]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111001100111111111101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][6]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[14][6]~DUPLICATE_q\,
	datad => \ALT_INV_RegFile[13][6]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux84~14_combout\,
	datag => \ALT_INV_RegFile[12][6]~q\,
	combout => \Mux84~1_combout\);

-- Location: LABCELL_X67_Y7_N6
\Mux84~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux84~13_combout\ = ( \Mux84~5_combout\ & ( \Mux84~1_combout\ & ( (!\R.curInst\(19) & (((\R.curInst\(18))) # (\Mux84~26_combout\))) # (\R.curInst\(19) & (((!\R.curInst\(18)) # (\Mux84~9_combout\)))) ) ) ) # ( !\Mux84~5_combout\ & ( \Mux84~1_combout\ & ( 
-- (!\R.curInst\(19) & (((\R.curInst\(18))) # (\Mux84~26_combout\))) # (\R.curInst\(19) & (((\Mux84~9_combout\ & \R.curInst\(18))))) ) ) ) # ( \Mux84~5_combout\ & ( !\Mux84~1_combout\ & ( (!\R.curInst\(19) & (\Mux84~26_combout\ & ((!\R.curInst\(18))))) # 
-- (\R.curInst\(19) & (((!\R.curInst\(18)) # (\Mux84~9_combout\)))) ) ) ) # ( !\Mux84~5_combout\ & ( !\Mux84~1_combout\ & ( (!\R.curInst\(19) & (\Mux84~26_combout\ & ((!\R.curInst\(18))))) # (\R.curInst\(19) & (((\Mux84~9_combout\ & \R.curInst\(18))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101000000000011010111110000001101010000111100110101111111110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux84~26_combout\,
	datab => \ALT_INV_Mux84~9_combout\,
	datac => \ALT_INV_R.curInst\(19),
	datad => \ALT_INV_R.curInst\(18),
	datae => \ALT_INV_Mux84~5_combout\,
	dataf => \ALT_INV_Mux84~1_combout\,
	combout => \Mux84~13_combout\);

-- Location: LABCELL_X73_Y7_N36
\Mux248~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux248~0_combout\ = ( \Mux84~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC\(6)))) ) ) # ( !\Mux84~13_combout\ & ( (\vAluSrc1~2_combout\ & (\R.curPC\(6) & !\vAluSrc1~1_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000000000000110000000011001111000000001100111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_vAluSrc1~2_combout\,
	datac => \ALT_INV_R.curPC\(6),
	datad => \ALT_INV_vAluSrc1~1_combout\,
	dataf => \ALT_INV_Mux84~13_combout\,
	combout => \Mux248~0_combout\);

-- Location: LABCELL_X74_Y7_N18
\ShiftLeft0~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~10_combout\ = ( \Mux247~0_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (\Mux248~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & ((\Mux249~0_combout\))) ) ) ) # ( !\Mux247~0_combout\ & ( 
-- \NxR.aluData2[1]~17_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (\Mux248~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & ((\Mux249~0_combout\))) ) ) ) # ( \Mux247~0_combout\ & ( !\NxR.aluData2[1]~17_combout\ & ( (\NxR.aluData2[0]~16_combout\) # 
-- (\Mux246~0_combout\) ) ) ) # ( !\Mux247~0_combout\ & ( !\NxR.aluData2[1]~17_combout\ & ( (\Mux246~0_combout\ & !\NxR.aluData2[0]~16_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100000000001100111111111101010101000011110101010100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux248~0_combout\,
	datab => \ALT_INV_Mux246~0_combout\,
	datac => \ALT_INV_Mux249~0_combout\,
	datad => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datae => \ALT_INV_Mux247~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[1]~17_combout\,
	combout => \ShiftLeft0~10_combout\);

-- Location: FF_X74_Y7_N19
\ShiftLeft0~10_NEW_REG210\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~10_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~10_OTERM211\);

-- Location: LABCELL_X81_Y8_N36
\ShiftLeft0~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~25_combout\ = ( \ShiftLeft0~24_OTERM293\ & ( \ShiftLeft0~5_OTERM203\ & ( (!\R.aluData2\(3) & (((!\R.aluData2\(2)) # (\ShiftLeft0~16_OTERM287\)))) # (\R.aluData2\(3) & (((\R.aluData2\(2))) # (\ShiftLeft0~10_OTERM211\))) ) ) ) # ( 
-- !\ShiftLeft0~24_OTERM293\ & ( \ShiftLeft0~5_OTERM203\ & ( (!\R.aluData2\(3) & (((\R.aluData2\(2) & \ShiftLeft0~16_OTERM287\)))) # (\R.aluData2\(3) & (((\R.aluData2\(2))) # (\ShiftLeft0~10_OTERM211\))) ) ) ) # ( \ShiftLeft0~24_OTERM293\ & ( 
-- !\ShiftLeft0~5_OTERM203\ & ( (!\R.aluData2\(3) & (((!\R.aluData2\(2)) # (\ShiftLeft0~16_OTERM287\)))) # (\R.aluData2\(3) & (\ShiftLeft0~10_OTERM211\ & (!\R.aluData2\(2)))) ) ) ) # ( !\ShiftLeft0~24_OTERM293\ & ( !\ShiftLeft0~5_OTERM203\ & ( 
-- (!\R.aluData2\(3) & (((\R.aluData2\(2) & \ShiftLeft0~16_OTERM287\)))) # (\R.aluData2\(3) & (\ShiftLeft0~10_OTERM211\ & (!\R.aluData2\(2)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000000011100110100001101110000010011000111111101001111011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~10_OTERM211\,
	datab => \ALT_INV_R.aluData2\(3),
	datac => \ALT_INV_R.aluData2\(2),
	datad => \ALT_INV_ShiftLeft0~16_OTERM287\,
	datae => \ALT_INV_ShiftLeft0~24_OTERM293\,
	dataf => \ALT_INV_ShiftLeft0~5_OTERM203\,
	combout => \ShiftLeft0~25_combout\);

-- Location: MLABCELL_X72_Y5_N6
\Selector16~1_RTM0795\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector16~1_RTM0795_combout\ = ( \Mux238~0_combout\ & ( ((!\NxR.aluData2[16]~5_combout\ & (\R.aluOp.ALUOpXor_OTERM355\)) # (\NxR.aluData2[16]~5_combout\ & ((\R.aluOp.ALUOpAnd_OTERM357\)))) # (\R.aluOp.ALUOpOr_OTERM353\) ) ) # ( !\Mux238~0_combout\ & ( 
-- (\NxR.aluData2[16]~5_combout\ & ((\R.aluOp.ALUOpXor_OTERM355\) # (\R.aluOp.ALUOpOr_OTERM353\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000011100000111000001110000011101110101011111110111010101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpOr_OTERM353\,
	datab => \ALT_INV_R.aluOp.ALUOpXor_OTERM355\,
	datac => \ALT_INV_NxR.aluData2[16]~5_combout\,
	datad => \ALT_INV_R.aluOp.ALUOpAnd_OTERM357\,
	dataf => \ALT_INV_Mux238~0_combout\,
	combout => \Selector16~1_RTM0795_combout\);

-- Location: FF_X72_Y5_N7
\Selector16~1_NEW_REG792\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector16~1_RTM0795_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector16~1_OTERM793\);

-- Location: LABCELL_X80_Y7_N36
\Selector16~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector16~2_combout\ = ( !\Selector17~0_OTERM391\ & ( \ShiftLeft0~0_OTERM263\ & ( (!\Selector16~1_OTERM793\ & !\Selector16~0_OTERM393\) ) ) ) # ( !\Selector17~0_OTERM391\ & ( !\ShiftLeft0~0_OTERM263\ & ( !\Selector16~1_OTERM793\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1100110011001100000000000000000011001100000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Selector16~1_OTERM793\,
	datad => \ALT_INV_Selector16~0_OTERM393\,
	datae => \ALT_INV_Selector17~0_OTERM391\,
	dataf => \ALT_INV_ShiftLeft0~0_OTERM263\,
	combout => \Selector16~2_combout\);

-- Location: LABCELL_X81_Y8_N24
\ShiftRight1~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~4_combout\ = ( \R.aluData2\(3) & ( \R.aluData2\(2) & ( \ShiftRight1~3_OTERM13\ ) ) ) # ( !\R.aluData2\(3) & ( \R.aluData2\(2) & ( \ShiftRight1~1_OTERM33\ ) ) ) # ( \R.aluData2\(3) & ( !\R.aluData2\(2) & ( \ShiftRight1~2_OTERM49\ ) ) ) # ( 
-- !\R.aluData2\(3) & ( !\R.aluData2\(2) & ( \ShiftRight1~0_OTERM257\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111010101010101010100000000111111110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~2_OTERM49\,
	datab => \ALT_INV_ShiftRight1~3_OTERM13\,
	datac => \ALT_INV_ShiftRight1~0_OTERM257\,
	datad => \ALT_INV_ShiftRight1~1_OTERM33\,
	datae => \ALT_INV_R.aluData2\(3),
	dataf => \ALT_INV_R.aluData2\(2),
	combout => \ShiftRight1~4_combout\);

-- Location: LABCELL_X81_Y8_N54
\Selector16~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector16~3_combout\ = ( \Selector16~2_combout\ & ( \ShiftRight1~4_combout\ & ( ((!\Selector31~0_OTERM349\ & ((!\ShiftLeft0~25_combout\) # (!\R.aluOp.ALUOpSLL~q\)))) # (\R.aluData2\(4)) ) ) ) # ( \Selector16~2_combout\ & ( !\ShiftRight1~4_combout\ & ( 
-- (!\ShiftLeft0~25_combout\) # ((!\R.aluOp.ALUOpSLL~q\) # (\R.aluData2\(4))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111010111100000000000000001100111110001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~25_combout\,
	datab => \ALT_INV_Selector31~0_OTERM349\,
	datac => \ALT_INV_R.aluData2\(4),
	datad => \ALT_INV_R.aluOp.ALUOpSLL~q\,
	datae => \ALT_INV_Selector16~2_combout\,
	dataf => \ALT_INV_ShiftRight1~4_combout\,
	combout => \Selector16~3_combout\);

-- Location: MLABCELL_X82_Y4_N0
\Selector16~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector16~5_combout\ = ( \Add1~65_sumout\ & ( \Add2~65_sumout\ & ( (!\Selector16~3_combout\) # ((\R.aluOp.ALUOpAdd~q\) # (\R.aluOp.ALUOpSub~q\)) ) ) ) # ( !\Add1~65_sumout\ & ( \Add2~65_sumout\ & ( (!\Selector16~3_combout\) # (\R.aluOp.ALUOpSub~q\) ) ) 
-- ) # ( \Add1~65_sumout\ & ( !\Add2~65_sumout\ & ( (!\Selector16~3_combout\) # (\R.aluOp.ALUOpAdd~q\) ) ) ) # ( !\Add1~65_sumout\ & ( !\Add2~65_sumout\ & ( !\Selector16~3_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010101010101010101011111010111110111011101110111011111110111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector16~3_combout\,
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datae => \ALT_INV_Add1~65_sumout\,
	dataf => \ALT_INV_Add2~65_sumout\,
	combout => \Selector16~5_combout\);

-- Location: LABCELL_X81_Y4_N6
\Comb:vJumpAdr[16]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[16]~0_combout\ = ( \R.aluRes\(16) & ( \Add3~65_sumout\ & ( (!\R.aluCalc~q\) # ((!\Equal4~2_combout\) # (\Selector16~5_combout\)) ) ) ) # ( !\R.aluRes\(16) & ( \Add3~65_sumout\ & ( (!\Equal4~2_combout\) # ((\R.aluCalc~q\ & 
-- \Selector16~5_combout\)) ) ) ) # ( \R.aluRes\(16) & ( !\Add3~65_sumout\ & ( (\Equal4~2_combout\ & ((!\R.aluCalc~q\) # (\Selector16~5_combout\))) ) ) ) # ( !\R.aluRes\(16) & ( !\Add3~65_sumout\ & ( (\R.aluCalc~q\ & (\Selector16~5_combout\ & 
-- \Equal4~2_combout\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000100000001000010110000101111110001111100011111101111111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluCalc~q\,
	datab => \ALT_INV_Selector16~5_combout\,
	datac => \ALT_INV_Equal4~2_combout\,
	datae => \ALT_INV_R.aluRes\(16),
	dataf => \ALT_INV_Add3~65_sumout\,
	combout => \Comb:vJumpAdr[16]~0_combout\);

-- Location: FF_X81_Y4_N8
\R.curPC[16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[16]~0_combout\,
	asdata => \Add0~57_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(16));

-- Location: FF_X63_Y3_N2
\RegFile[14][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][16]~q\);

-- Location: LABCELL_X63_Y1_N12
\Mux74~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux74~14_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[8][16]~q\))) # (\R.curInst\(15) & (\RegFile[9][16]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & (\RegFile[10][16]~q\)) # (\R.curInst\(15) & ((\RegFile[11][16]~q\))))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][16]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[10][16]~q\,
	datad => \ALT_INV_RegFile[11][16]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][16]~q\,
	combout => \Mux74~14_combout\);

-- Location: FF_X63_Y3_N23
\RegFile[12][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][16]~q\);

-- Location: LABCELL_X63_Y3_N12
\Mux74~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux74~1_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux74~14_combout\)))) # (\R.curInst\(17) & ((!\Mux74~14_combout\ & ((\RegFile[12][16]~q\))) # (\Mux74~14_combout\ & (\RegFile[13][16]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux74~14_combout\)))) # (\R.curInst\(17) & ((!\Mux74~14_combout\ & ((\RegFile[14][16]~q\))) # (\Mux74~14_combout\ & (\RegFile[15][16]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][16]~q\,
	datab => \ALT_INV_RegFile[15][16]~q\,
	datac => \ALT_INV_RegFile[14][16]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux74~14_combout\,
	datag => \ALT_INV_RegFile[12][16]~q\,
	combout => \Mux74~1_combout\);

-- Location: MLABCELL_X65_Y2_N18
\Mux74~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux74~18_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & (\RegFile[16][16]~q\)) # (\R.curInst\(15) & ((\RegFile[17][16]~q\)))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & ((\RegFile[18][16]~q\))) # (\R.curInst\(15) & (\RegFile[19][16]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001010101111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[19][16]~q\,
	datac => \ALT_INV_RegFile[18][16]~q\,
	datad => \ALT_INV_RegFile[17][16]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][16]~q\,
	combout => \Mux74~18_combout\);

-- Location: FF_X71_Y1_N55
\RegFile[20][16]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][16]~DUPLICATE_q\);

-- Location: MLABCELL_X65_Y2_N54
\Mux74~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux74~5_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux74~18_combout\)))) # (\R.curInst\(17) & ((!\Mux74~18_combout\ & ((\RegFile[20][16]~DUPLICATE_q\))) # (\Mux74~18_combout\ & (\RegFile[21][16]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux74~18_combout\)))) # (\R.curInst\(17) & ((!\Mux74~18_combout\ & ((\RegFile[22][16]~q\))) # (\Mux74~18_combout\ & (\RegFile[23][16]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[23][16]~q\,
	datab => \ALT_INV_RegFile[21][16]~q\,
	datac => \ALT_INV_RegFile[22][16]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux74~18_combout\,
	datag => \ALT_INV_RegFile[20][16]~DUPLICATE_q\,
	combout => \Mux74~5_combout\);

-- Location: FF_X68_Y3_N11
\RegFile[5][16]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(16),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][16]~q\);

-- Location: LABCELL_X68_Y3_N48
\Mux74~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux74~0_combout\ = ( \RegFile[7][16]~q\ & ( \R.curInst\(15) & ( (\RegFile[5][16]~q\) # (\R.curInst\(16)) ) ) ) # ( !\RegFile[7][16]~q\ & ( \R.curInst\(15) & ( (!\R.curInst\(16) & \RegFile[5][16]~q\) ) ) ) # ( \RegFile[7][16]~q\ & ( !\R.curInst\(15) & ( 
-- (!\R.curInst\(16) & (\RegFile[4][16]~q\)) # (\R.curInst\(16) & ((\RegFile[6][16]~q\))) ) ) ) # ( !\RegFile[7][16]~q\ & ( !\R.curInst\(15) & ( (!\R.curInst\(16) & (\RegFile[4][16]~q\)) # (\R.curInst\(16) & ((\RegFile[6][16]~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101001101010011010100110101001100000000111100000000111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[4][16]~q\,
	datab => \ALT_INV_RegFile[6][16]~q\,
	datac => \ALT_INV_R.curInst\(16),
	datad => \ALT_INV_RegFile[5][16]~q\,
	datae => \ALT_INV_RegFile[7][16]~q\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux74~0_combout\);

-- Location: LABCELL_X68_Y3_N42
\Mux74~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux74~26_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (\R.curInst\(15) & (\RegFile[1][16]~q\))) # (\R.curInst\(17) & ((((\Mux74~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & ((!\R.curInst\(15) & (\RegFile[2][16]~q\)) # 
-- (\R.curInst\(15) & (((\RegFile[3][16]~q\)))))) # (\R.curInst\(17) & ((((\Mux74~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001000000010000010000010101001010111010101110101110101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_R.curInst\(15),
	datac => \ALT_INV_RegFile[2][16]~q\,
	datad => \ALT_INV_RegFile[3][16]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux74~0_combout\,
	datag => \ALT_INV_RegFile[1][16]~q\,
	combout => \Mux74~26_combout\);

-- Location: LABCELL_X66_Y2_N12
\Mux74~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux74~22_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[24][16]~q\))) # (\R.curInst\(15) & (\RegFile[25][16]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[26][16]~q\))) # (\R.curInst\(15) & (\RegFile[27][16]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[25][16]~q\,
	datab => \ALT_INV_RegFile[27][16]~q\,
	datac => \ALT_INV_RegFile[26][16]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][16]~q\,
	combout => \Mux74~22_combout\);

-- Location: LABCELL_X67_Y5_N0
\Mux74~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux74~9_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux74~22_combout\)))) # (\R.curInst\(17) & ((!\Mux74~22_combout\ & ((\RegFile[28][16]~q\))) # (\Mux74~22_combout\ & (\RegFile[29][16]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux74~22_combout\)))) # (\R.curInst\(17) & ((!\Mux74~22_combout\ & ((\RegFile[30][16]~q\))) # (\Mux74~22_combout\ & (\RegFile[31][16]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][16]~q\,
	datab => \ALT_INV_RegFile[29][16]~q\,
	datac => \ALT_INV_RegFile[30][16]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux74~22_combout\,
	datag => \ALT_INV_RegFile[28][16]~q\,
	combout => \Mux74~9_combout\);

-- Location: LABCELL_X67_Y3_N45
\Mux74~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux74~13_combout\ = ( \Mux74~26_combout\ & ( \Mux74~9_combout\ & ( (!\R.curInst\(18) & ((!\R.curInst\(19)) # ((\Mux74~5_combout\)))) # (\R.curInst\(18) & (((\Mux74~1_combout\)) # (\R.curInst\(19)))) ) ) ) # ( !\Mux74~26_combout\ & ( \Mux74~9_combout\ & ( 
-- (!\R.curInst\(18) & (\R.curInst\(19) & ((\Mux74~5_combout\)))) # (\R.curInst\(18) & (((\Mux74~1_combout\)) # (\R.curInst\(19)))) ) ) ) # ( \Mux74~26_combout\ & ( !\Mux74~9_combout\ & ( (!\R.curInst\(18) & ((!\R.curInst\(19)) # ((\Mux74~5_combout\)))) # 
-- (\R.curInst\(18) & (!\R.curInst\(19) & (\Mux74~1_combout\))) ) ) ) # ( !\Mux74~26_combout\ & ( !\Mux74~9_combout\ & ( (!\R.curInst\(18) & (\R.curInst\(19) & ((\Mux74~5_combout\)))) # (\R.curInst\(18) & (!\R.curInst\(19) & (\Mux74~1_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010000100110100011001010111000010101001101111001110110111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(18),
	datab => \ALT_INV_R.curInst\(19),
	datac => \ALT_INV_Mux74~1_combout\,
	datad => \ALT_INV_Mux74~5_combout\,
	datae => \ALT_INV_Mux74~26_combout\,
	dataf => \ALT_INV_Mux74~9_combout\,
	combout => \Mux74~13_combout\);

-- Location: LABCELL_X73_Y6_N3
\Mux238~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux238~0_combout\ = ( \Mux74~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC\(16)))) ) ) # ( !\Mux74~13_combout\ & ( (\vAluSrc1~2_combout\ & (!\vAluSrc1~1_combout\ & \R.curPC\(16))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110000000000000011000011000000111100001100000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_vAluSrc1~2_combout\,
	datac => \ALT_INV_vAluSrc1~1_combout\,
	datad => \ALT_INV_R.curPC\(16),
	dataf => \ALT_INV_Mux74~13_combout\,
	combout => \Mux238~0_combout\);

-- Location: LABCELL_X73_Y6_N30
\ShiftRight1~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~18_combout\ = ( \Mux239~0_combout\ & ( \Mux240~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((\Mux241~0_combout\) # (\NxR.aluData2[0]~16_combout\)))) # (\NxR.aluData2[1]~17_combout\ & (((!\NxR.aluData2[0]~16_combout\)) # 
-- (\Mux238~0_combout\))) ) ) ) # ( !\Mux239~0_combout\ & ( \Mux240~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((\Mux241~0_combout\) # (\NxR.aluData2[0]~16_combout\)))) # (\NxR.aluData2[1]~17_combout\ & (\Mux238~0_combout\ & 
-- (\NxR.aluData2[0]~16_combout\))) ) ) ) # ( \Mux239~0_combout\ & ( !\Mux240~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((!\NxR.aluData2[0]~16_combout\ & \Mux241~0_combout\)))) # (\NxR.aluData2[1]~17_combout\ & (((!\NxR.aluData2[0]~16_combout\)) # 
-- (\Mux238~0_combout\))) ) ) ) # ( !\Mux239~0_combout\ & ( !\Mux240~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (((!\NxR.aluData2[0]~16_combout\ & \Mux241~0_combout\)))) # (\NxR.aluData2[1]~17_combout\ & (\Mux238~0_combout\ & 
-- (\NxR.aluData2[0]~16_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000111000001001100011111000100001101110011010011110111111101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux238~0_combout\,
	datab => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datac => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datad => \ALT_INV_Mux241~0_combout\,
	datae => \ALT_INV_Mux239~0_combout\,
	dataf => \ALT_INV_Mux240~0_combout\,
	combout => \ShiftRight1~18_combout\);

-- Location: FF_X73_Y6_N31
\ShiftRight1~18_NEW_REG268\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~18_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~18_OTERM269\);

-- Location: MLABCELL_X78_Y9_N18
\ShiftRight1~47\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~47_combout\ = ( \ShiftRight1~17_OTERM267\ & ( \ShiftRight1~10_OTERM265\ & ( (!\R.aluData2\(2)) # ((!\R.aluData2\(3) & (\ShiftRight1~18_OTERM269\)) # (\R.aluData2\(3) & ((\ShiftRight1~11_OTERM35\)))) ) ) ) # ( !\ShiftRight1~17_OTERM267\ & ( 
-- \ShiftRight1~10_OTERM265\ & ( (!\R.aluData2\(3) & (\ShiftRight1~18_OTERM269\ & ((\R.aluData2\(2))))) # (\R.aluData2\(3) & (((!\R.aluData2\(2)) # (\ShiftRight1~11_OTERM35\)))) ) ) ) # ( \ShiftRight1~17_OTERM267\ & ( !\ShiftRight1~10_OTERM265\ & ( 
-- (!\R.aluData2\(3) & (((!\R.aluData2\(2))) # (\ShiftRight1~18_OTERM269\))) # (\R.aluData2\(3) & (((\ShiftRight1~11_OTERM35\ & \R.aluData2\(2))))) ) ) ) # ( !\ShiftRight1~17_OTERM267\ & ( !\ShiftRight1~10_OTERM265\ & ( (\R.aluData2\(2) & ((!\R.aluData2\(3) 
-- & (\ShiftRight1~18_OTERM269\)) # (\R.aluData2\(3) & ((\ShiftRight1~11_OTERM35\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001000111110011000100011100110011010001111111111101000111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~18_OTERM269\,
	datab => \ALT_INV_R.aluData2\(3),
	datac => \ALT_INV_ShiftRight1~11_OTERM35\,
	datad => \ALT_INV_R.aluData2\(2),
	datae => \ALT_INV_ShiftRight1~17_OTERM267\,
	dataf => \ALT_INV_ShiftRight1~10_OTERM265\,
	combout => \ShiftRight1~47_combout\);

-- Location: LABCELL_X79_Y9_N3
\Selector23~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector23~5_combout\ = ( \Selector23~4_combout\ & ( !\Selector23~2_combout\ & ( (!\Selector23~1_combout\ & ((!\Selector31~5_OTERM599\) # (!\ShiftRight1~47_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111000001110000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector31~5_OTERM599\,
	datab => \ALT_INV_ShiftRight1~47_combout\,
	datac => \ALT_INV_Selector23~1_combout\,
	datae => \ALT_INV_Selector23~4_combout\,
	dataf => \ALT_INV_Selector23~2_combout\,
	combout => \Selector23~5_combout\);

-- Location: LABCELL_X80_Y3_N24
\Selector23~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector23~0_combout\ = ( \Add1~37_sumout\ & ( ((\R.aluOp.ALUOpSub~q\ & \Add2~37_sumout\)) # (\R.aluOp.ALUOpAdd~q\) ) ) # ( !\Add1~37_sumout\ & ( (\R.aluOp.ALUOpSub~q\ & \Add2~37_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101000001010000010100110111001101110011011100110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datab => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datac => \ALT_INV_Add2~37_sumout\,
	dataf => \ALT_INV_Add1~37_sumout\,
	combout => \Selector23~0_combout\);

-- Location: LABCELL_X77_Y3_N42
\Comb:vJumpAdr[9]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[9]~0_combout\ = ( \Equal4~2_combout\ & ( \Add3~37_sumout\ & ( (!\R.aluCalc~q\ & (((\R.aluRes\(9))))) # (\R.aluCalc~q\ & ((!\Selector23~5_combout\) # ((\Selector23~0_combout\)))) ) ) ) # ( !\Equal4~2_combout\ & ( \Add3~37_sumout\ ) ) # ( 
-- \Equal4~2_combout\ & ( !\Add3~37_sumout\ & ( (!\R.aluCalc~q\ & (((\R.aluRes\(9))))) # (\R.aluCalc~q\ & ((!\Selector23~5_combout\) # ((\Selector23~0_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000001110100011111111111111111111110011101000111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector23~5_combout\,
	datab => \ALT_INV_R.aluRes\(9),
	datac => \ALT_INV_R.aluCalc~q\,
	datad => \ALT_INV_Selector23~0_combout\,
	datae => \ALT_INV_Equal4~2_combout\,
	dataf => \ALT_INV_Add3~37_sumout\,
	combout => \Comb:vJumpAdr[9]~0_combout\);

-- Location: FF_X77_Y3_N43
\R.curPC[9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[9]~0_combout\,
	asdata => \Add0~29_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(9));

-- Location: LABCELL_X81_Y6_N24
\Add0~33\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~33_sumout\ = SUM(( \R.curPC\(10) ) + ( GND ) + ( \Add0~30\ ))
-- \Add0~34\ = CARRY(( \R.curPC\(10) ) + ( GND ) + ( \Add0~30\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.curPC\(10),
	cin => \Add0~30\,
	sumout => \Add0~33_sumout\,
	cout => \Add0~34\);

-- Location: LABCELL_X80_Y8_N18
\R.regWriteData[10]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.regWriteData[10]~feeder_combout\ = \Add0~33_sumout\

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110011001100110011001100110011001100110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Add0~33_sumout\,
	combout => \R.regWriteData[10]~feeder_combout\);

-- Location: MLABCELL_X82_Y6_N48
\ShiftRight1~49\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~49_combout\ = ( \ShiftRight1~22_OTERM273\ & ( \ShiftRight1~25_OTERM277\ & ( (!\R.aluData2\(2)) # ((!\R.aluData2\(3) & ((\ShiftRight1~23_OTERM275\))) # (\R.aluData2\(3) & (\ShiftRight1~26_OTERM37\))) ) ) ) # ( !\ShiftRight1~22_OTERM273\ & ( 
-- \ShiftRight1~25_OTERM277\ & ( (!\R.aluData2\(3) & (((\R.aluData2\(2) & \ShiftRight1~23_OTERM275\)))) # (\R.aluData2\(3) & (((!\R.aluData2\(2))) # (\ShiftRight1~26_OTERM37\))) ) ) ) # ( \ShiftRight1~22_OTERM273\ & ( !\ShiftRight1~25_OTERM277\ & ( 
-- (!\R.aluData2\(3) & (((!\R.aluData2\(2)) # (\ShiftRight1~23_OTERM275\)))) # (\R.aluData2\(3) & (\ShiftRight1~26_OTERM37\ & (\R.aluData2\(2)))) ) ) ) # ( !\ShiftRight1~22_OTERM273\ & ( !\ShiftRight1~25_OTERM277\ & ( (\R.aluData2\(2) & ((!\R.aluData2\(3) & 
-- ((\ShiftRight1~23_OTERM275\))) # (\R.aluData2\(3) & (\ShiftRight1~26_OTERM37\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000100001101110000011100110100110001001111011111000111111101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~26_OTERM37\,
	datab => \ALT_INV_R.aluData2\(3),
	datac => \ALT_INV_R.aluData2\(2),
	datad => \ALT_INV_ShiftRight1~23_OTERM275\,
	datae => \ALT_INV_ShiftRight1~22_OTERM273\,
	dataf => \ALT_INV_ShiftRight1~25_OTERM277\,
	combout => \ShiftRight1~49_combout\);

-- Location: LABCELL_X77_Y8_N36
\Selector22~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector22~3_combout\ = ( \R.aluData2\(2) & ( \R.aluOp.ALUOpSLL~q\ & ( (\ShiftLeft0~8_OTERM207\ & !\R.aluData2\(3)) ) ) ) # ( !\R.aluData2\(2) & ( \R.aluOp.ALUOpSLL~q\ & ( (!\R.aluData2\(3) & ((\ShiftLeft0~13_OTERM285\))) # (\R.aluData2\(3) & 
-- (\ShiftLeft0~2_OTERM221\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000011110011110100010001000100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~8_OTERM207\,
	datab => \ALT_INV_R.aluData2\(3),
	datac => \ALT_INV_ShiftLeft0~2_OTERM221\,
	datad => \ALT_INV_ShiftLeft0~13_OTERM285\,
	datae => \ALT_INV_R.aluData2\(2),
	dataf => \ALT_INV_R.aluOp.ALUOpSLL~q\,
	combout => \Selector22~3_combout\);

-- Location: LABCELL_X80_Y8_N42
\Selector22~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector22~4_combout\ = ( \Selector31~0_OTERM349\ & ( \Add1~41_sumout\ & ( ((!\R.aluData2\(4) & ((\Selector22~3_combout\) # (\ShiftRight1~49_combout\)))) # (\R.aluOp.ALUOpAdd~q\) ) ) ) # ( !\Selector31~0_OTERM349\ & ( \Add1~41_sumout\ & ( 
-- ((\Selector22~3_combout\ & !\R.aluData2\(4))) # (\R.aluOp.ALUOpAdd~q\) ) ) ) # ( \Selector31~0_OTERM349\ & ( !\Add1~41_sumout\ & ( (!\R.aluData2\(4) & ((\Selector22~3_combout\) # (\ShiftRight1~49_combout\))) ) ) ) # ( !\Selector31~0_OTERM349\ & ( 
-- !\Add1~41_sumout\ & ( (\Selector22~3_combout\ & !\R.aluData2\(4)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100000000010111110000000000111111001100110111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~49_combout\,
	datab => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datac => \ALT_INV_Selector22~3_combout\,
	datad => \ALT_INV_R.aluData2\(4),
	datae => \ALT_INV_Selector31~0_OTERM349\,
	dataf => \ALT_INV_Add1~41_sumout\,
	combout => \Selector22~4_combout\);

-- Location: LABCELL_X80_Y8_N12
\Selector22~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector22~2_combout\ = ( \Selector22~0_RTM0477_combout\ & ( \Add2~41_sumout\ & ( (!\R.aluOp.ALUOpSub~q\ & (!\Selector22~1_OTERM427\ & !\R.aluData2\(4))) ) ) ) # ( !\Selector22~0_RTM0477_combout\ & ( \Add2~41_sumout\ & ( (!\R.aluOp.ALUOpSub~q\ & 
-- !\Selector22~1_OTERM427\) ) ) ) # ( \Selector22~0_RTM0477_combout\ & ( !\Add2~41_sumout\ & ( (!\Selector22~1_OTERM427\ & !\R.aluData2\(4)) ) ) ) # ( !\Selector22~0_RTM0477_combout\ & ( !\Add2~41_sumout\ & ( !\Selector22~1_OTERM427\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111000011110000111100000000000011000000110000001100000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_Selector22~1_OTERM427\,
	datad => \ALT_INV_R.aluData2\(4),
	datae => \ALT_INV_Selector22~0_RTM0477_combout\,
	dataf => \ALT_INV_Add2~41_sumout\,
	combout => \Selector22~2_combout\);

-- Location: LABCELL_X81_Y8_N18
\Selector22~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector22~5_combout\ = ( \Selector22~2_combout\ & ( \Selector22~4_combout\ ) ) # ( !\Selector22~2_combout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111001100110011001111111111111111110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Selector22~4_combout\,
	datae => \ALT_INV_Selector22~2_combout\,
	combout => \Selector22~5_combout\);

-- Location: FF_X81_Y8_N19
\R.aluRes[10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector22~5_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(10));

-- Location: IOIBUF_X56_Y0_N52
\avm_d_readdata[18]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(18),
	o => \avm_d_readdata[18]~input_o\);

-- Location: LABCELL_X79_Y2_N12
\Comb:vRegWriteData[10]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[10]~0_combout\ = ( !\R.curInst\(13) & ( \R.curInst\(12) & ( \avm_d_readdata[18]~input_o\ ) ) ) # ( \R.curInst\(13) & ( !\R.curInst\(12) & ( (!\R.curInst\(14) & \avm_d_readdata[18]~input_o\) ) ) ) # ( !\R.curInst\(13) & ( 
-- !\R.curInst\(12) & ( (!\R.curInst\(14) & \avm_d_readdata[31]~input_o\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010001000100010000010100000101000001111000011110000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(14),
	datab => \ALT_INV_avm_d_readdata[31]~input_o\,
	datac => \ALT_INV_avm_d_readdata[18]~input_o\,
	datae => \ALT_INV_R.curInst\(13),
	dataf => \ALT_INV_R.curInst\(12),
	combout => \Comb:vRegWriteData[10]~0_combout\);

-- Location: LABCELL_X80_Y8_N54
\Comb:vRegWriteData[10]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[10]~1_combout\ = ( \R.aluCalc~q\ & ( \Comb:vRegWriteData[10]~0_combout\ & ( (!\Selector22~2_combout\) # ((\Selector22~4_combout\) # (\R.memToReg~q\)) ) ) ) # ( !\R.aluCalc~q\ & ( \Comb:vRegWriteData[10]~0_combout\ & ( (\R.memToReg~q\) 
-- # (\R.aluRes\(10)) ) ) ) # ( \R.aluCalc~q\ & ( !\Comb:vRegWriteData[10]~0_combout\ & ( (!\R.memToReg~q\ & ((!\Selector22~2_combout\) # (\Selector22~4_combout\))) ) ) ) # ( !\R.aluCalc~q\ & ( !\Comb:vRegWriteData[10]~0_combout\ & ( (\R.aluRes\(10) & 
-- !\R.memToReg~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101000001010000110000001111000001011111010111111100111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluRes\(10),
	datab => \ALT_INV_Selector22~2_combout\,
	datac => \ALT_INV_R.memToReg~q\,
	datad => \ALT_INV_Selector22~4_combout\,
	datae => \ALT_INV_R.aluCalc~q\,
	dataf => \ALT_INV_Comb:vRegWriteData[10]~0_combout\,
	combout => \Comb:vRegWriteData[10]~1_combout\);

-- Location: FF_X80_Y8_N20
\R.regWriteData[10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \R.regWriteData[10]~feeder_combout\,
	asdata => \Comb:vRegWriteData[10]~1_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(10));

-- Location: FF_X65_Y6_N8
\RegFile[2][10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(10),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][10]~q\);

-- Location: MLABCELL_X65_Y6_N24
\Mux112~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux112~0_combout\ = ( \RegFile[6][10]~q\ & ( \R.curInst\(21) & ( (!\R.curInst\(20)) # (\RegFile[7][10]~q\) ) ) ) # ( !\RegFile[6][10]~q\ & ( \R.curInst\(21) & ( (\R.curInst\(20) & \RegFile[7][10]~q\) ) ) ) # ( \RegFile[6][10]~q\ & ( !\R.curInst\(21) & ( 
-- (!\R.curInst\(20) & (\RegFile[4][10]~q\)) # (\R.curInst\(20) & ((\RegFile[5][10]~q\))) ) ) ) # ( !\RegFile[6][10]~q\ & ( !\R.curInst\(21) & ( (!\R.curInst\(20) & (\RegFile[4][10]~q\)) # (\R.curInst\(20) & ((\RegFile[5][10]~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101001011111000010100101111100010001000100011011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(20),
	datab => \ALT_INV_RegFile[7][10]~q\,
	datac => \ALT_INV_RegFile[4][10]~q\,
	datad => \ALT_INV_RegFile[5][10]~q\,
	datae => \ALT_INV_RegFile[6][10]~q\,
	dataf => \ALT_INV_R.curInst\(21),
	combout => \Mux112~0_combout\);

-- Location: MLABCELL_X65_Y6_N6
\Mux112~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux112~26_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (\R.curInst\(20) & (\RegFile[1][10]~q\))) # (\R.curInst\(22) & ((((\Mux112~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (\RegFile[2][10]~q\)) # 
-- (\R.curInst\(20) & (((\RegFile[3][10]~q\)))))) # (\R.curInst\(22) & ((((\Mux112~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010000000100000010000100110000110111001101110011101101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(20),
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[2][10]~q\,
	datad => \ALT_INV_RegFile[3][10]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux112~0_combout\,
	datag => \ALT_INV_RegFile[1][10]~q\,
	combout => \Mux112~26_combout\);

-- Location: LABCELL_X66_Y6_N12
\Mux112~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux112~22_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[24][10]~q\))) # (\R.curInst\(20) & (\RegFile[25][10]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[26][10]~q\))) # (\R.curInst\(20) & (\RegFile[27][10]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[25][10]~q\,
	datab => \ALT_INV_RegFile[27][10]~q\,
	datac => \ALT_INV_RegFile[26][10]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][10]~q\,
	combout => \Mux112~22_combout\);

-- Location: LABCELL_X66_Y6_N54
\Mux112~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux112~9_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux112~22_combout\)))) # (\R.curInst\(22) & ((!\Mux112~22_combout\ & ((\RegFile[28][10]~q\))) # (\Mux112~22_combout\ & (\RegFile[29][10]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux112~22_combout\)))) # (\R.curInst\(22) & ((!\Mux112~22_combout\ & ((\RegFile[30][10]~q\))) # (\Mux112~22_combout\ & (\RegFile[31][10]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[29][10]~q\,
	datab => \ALT_INV_RegFile[31][10]~q\,
	datac => \ALT_INV_RegFile[30][10]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux112~22_combout\,
	datag => \ALT_INV_RegFile[28][10]~q\,
	combout => \Mux112~9_combout\);

-- Location: MLABCELL_X65_Y8_N24
\Mux112~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux112~18_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[16][10]~q\))) # (\R.curInst\(20) & (\RegFile[17][10]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[18][10]~q\))) # (\R.curInst\(20) & (\RegFile[19][10]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[19][10]~q\,
	datab => \ALT_INV_RegFile[17][10]~q\,
	datac => \ALT_INV_RegFile[18][10]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][10]~q\,
	combout => \Mux112~18_combout\);

-- Location: MLABCELL_X65_Y8_N30
\Mux112~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux112~5_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux112~18_combout\)))) # (\R.curInst\(22) & ((!\Mux112~18_combout\ & ((\RegFile[20][10]~q\))) # (\Mux112~18_combout\ & (\RegFile[21][10]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux112~18_combout\)))) # (\R.curInst\(22) & ((!\Mux112~18_combout\ & ((\RegFile[22][10]~q\))) # (\Mux112~18_combout\ & (\RegFile[23][10]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][10]~q\,
	datab => \ALT_INV_RegFile[23][10]~q\,
	datac => \ALT_INV_RegFile[22][10]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux112~18_combout\,
	datag => \ALT_INV_RegFile[20][10]~q\,
	combout => \Mux112~5_combout\);

-- Location: FF_X60_Y8_N37
\RegFile[10][10]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[10][10]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][10]~DUPLICATE_q\);

-- Location: LABCELL_X66_Y8_N33
\Mux112~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux112~14_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & (\RegFile[8][10]~q\)) # (\R.curInst\(20) & ((\RegFile[9][10]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & ((\RegFile[10][10]~DUPLICATE_q\))) # (\R.curInst\(20) & (\RegFile[11][10]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110000110011111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[11][10]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[10][10]~DUPLICATE_q\,
	datad => \ALT_INV_RegFile[9][10]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][10]~q\,
	combout => \Mux112~14_combout\);

-- Location: FF_X70_Y8_N1
\RegFile[12][10]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[12][10]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][10]~DUPLICATE_q\);

-- Location: LABCELL_X66_Y8_N18
\Mux112~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux112~1_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux112~14_combout\)))) # (\R.curInst\(22) & ((!\Mux112~14_combout\ & (\RegFile[12][10]~DUPLICATE_q\)) # (\Mux112~14_combout\ & ((\RegFile[13][10]~q\)))))) ) ) # ( \R.curInst\(21) & ( 
-- (!\R.curInst\(22) & ((((\Mux112~14_combout\))))) # (\R.curInst\(22) & (((!\Mux112~14_combout\ & ((\RegFile[14][10]~q\))) # (\Mux112~14_combout\ & (\RegFile[15][10]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111001100111111111101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][10]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[14][10]~q\,
	datad => \ALT_INV_RegFile[13][10]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux112~14_combout\,
	datag => \ALT_INV_RegFile[12][10]~DUPLICATE_q\,
	combout => \Mux112~1_combout\);

-- Location: LABCELL_X66_Y6_N36
\Mux112~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux112~13_combout\ = ( \Mux112~5_combout\ & ( \Mux112~1_combout\ & ( (!\R.curInst\(23) & (((\Mux112~26_combout\)) # (\R.curInst\(24)))) # (\R.curInst\(23) & ((!\R.curInst\(24)) # ((\Mux112~9_combout\)))) ) ) ) # ( !\Mux112~5_combout\ & ( 
-- \Mux112~1_combout\ & ( (!\R.curInst\(23) & (!\R.curInst\(24) & (\Mux112~26_combout\))) # (\R.curInst\(23) & ((!\R.curInst\(24)) # ((\Mux112~9_combout\)))) ) ) ) # ( \Mux112~5_combout\ & ( !\Mux112~1_combout\ & ( (!\R.curInst\(23) & 
-- (((\Mux112~26_combout\)) # (\R.curInst\(24)))) # (\R.curInst\(23) & (\R.curInst\(24) & ((\Mux112~9_combout\)))) ) ) ) # ( !\Mux112~5_combout\ & ( !\Mux112~1_combout\ & ( (!\R.curInst\(23) & (!\R.curInst\(24) & (\Mux112~26_combout\))) # (\R.curInst\(23) & 
-- (\R.curInst\(24) & ((\Mux112~9_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000100000011001001010100011101101001100010111010110111001111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(23),
	datab => \ALT_INV_R.curInst\(24),
	datac => \ALT_INV_Mux112~26_combout\,
	datad => \ALT_INV_Mux112~9_combout\,
	datae => \ALT_INV_Mux112~5_combout\,
	dataf => \ALT_INV_Mux112~1_combout\,
	combout => \Mux112~13_combout\);

-- Location: LABCELL_X75_Y6_N0
\NxR.aluData2[10]~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[10]~9_combout\ = ( \Mux112~13_combout\ & ( (!\vAluSrc2~1_combout\) # ((\Equal4~1_combout\ & \Mux144~0_combout\)) ) ) # ( !\Mux112~13_combout\ & ( (\Equal4~1_combout\ & (\Mux144~0_combout\ & \vAluSrc2~1_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000101000000000000010111111111000001011111111100000101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Equal4~1_combout\,
	datac => \ALT_INV_Mux144~0_combout\,
	datad => \ALT_INV_vAluSrc2~1_combout\,
	dataf => \ALT_INV_Mux112~13_combout\,
	combout => \NxR.aluData2[10]~9_combout\);

-- Location: LABCELL_X75_Y6_N57
\Selector22~1_RTM0429\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector22~1_RTM0429_combout\ = ( \Mux244~0_combout\ & ( ((!\NxR.aluData2[10]~9_combout\ & ((\R.aluOp.ALUOpXor_OTERM355\))) # (\NxR.aluData2[10]~9_combout\ & (\R.aluOp.ALUOpAnd_OTERM357\))) # (\R.aluOp.ALUOpOr_OTERM353\) ) ) # ( !\Mux244~0_combout\ & ( 
-- (\NxR.aluData2[10]~9_combout\ & ((\R.aluOp.ALUOpOr_OTERM353\) # (\R.aluOp.ALUOpXor_OTERM355\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000111111000000000011111100111111010111110011111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpAnd_OTERM357\,
	datab => \ALT_INV_R.aluOp.ALUOpXor_OTERM355\,
	datac => \ALT_INV_R.aluOp.ALUOpOr_OTERM353\,
	datad => \ALT_INV_NxR.aluData2[10]~9_combout\,
	dataf => \ALT_INV_Mux244~0_combout\,
	combout => \Selector22~1_RTM0429_combout\);

-- Location: FF_X75_Y6_N58
\Selector22~1_NEW_REG426\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector22~1_RTM0429_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector22~1_OTERM427\);

-- Location: LABCELL_X81_Y9_N39
\vAluRes~32\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~32_combout\ = ( \R.aluData2\(4) & ( \Selector22~0_RTM0477_combout\ & ( (\R.aluCalc~q\) # (\R.aluRes\(10)) ) ) ) # ( !\R.aluData2\(4) & ( \Selector22~0_RTM0477_combout\ & ( (\R.aluRes\(10) & !\R.aluCalc~q\) ) ) ) # ( \R.aluData2\(4) & ( 
-- !\Selector22~0_RTM0477_combout\ & ( (\R.aluRes\(10) & !\R.aluCalc~q\) ) ) ) # ( !\R.aluData2\(4) & ( !\Selector22~0_RTM0477_combout\ & ( (\R.aluRes\(10) & !\R.aluCalc~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011000000110000001100000011000000110000001100000011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluRes\(10),
	datac => \ALT_INV_R.aluCalc~q\,
	datae => \ALT_INV_R.aluData2\(4),
	dataf => \ALT_INV_Selector22~0_RTM0477_combout\,
	combout => \vAluRes~32_combout\);

-- Location: LABCELL_X80_Y8_N48
\vAluRes~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~10_combout\ = ( \R.aluOp.ALUOpSub~q\ & ( \Selector22~4_combout\ & ( (\R.aluCalc~q\) # (\vAluRes~32_combout\) ) ) ) # ( !\R.aluOp.ALUOpSub~q\ & ( \Selector22~4_combout\ & ( (\R.aluCalc~q\) # (\vAluRes~32_combout\) ) ) ) # ( \R.aluOp.ALUOpSub~q\ & 
-- ( !\Selector22~4_combout\ & ( ((\R.aluCalc~q\ & ((\Add2~41_sumout\) # (\Selector22~1_OTERM427\)))) # (\vAluRes~32_combout\) ) ) ) # ( !\R.aluOp.ALUOpSub~q\ & ( !\Selector22~4_combout\ & ( ((\Selector22~1_OTERM427\ & \R.aluCalc~q\)) # 
-- (\vAluRes~32_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001101110111001100110111111100110011111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector22~1_OTERM427\,
	datab => \ALT_INV_vAluRes~32_combout\,
	datac => \ALT_INV_Add2~41_sumout\,
	datad => \ALT_INV_R.aluCalc~q\,
	datae => \ALT_INV_R.aluOp.ALUOpSub~q\,
	dataf => \ALT_INV_Selector22~4_combout\,
	combout => \vAluRes~10_combout\);

-- Location: LABCELL_X80_Y8_N0
\Comb:vJumpAdr[10]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[10]~0_combout\ = ( \Add3~41_sumout\ & ( (!\Equal4~2_combout\) # (\vAluRes~10_combout\) ) ) # ( !\Add3~41_sumout\ & ( (\Equal4~2_combout\ & \vAluRes~10_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000110000001111001111110011111100111111001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Equal4~2_combout\,
	datac => \ALT_INV_vAluRes~10_combout\,
	dataf => \ALT_INV_Add3~41_sumout\,
	combout => \Comb:vJumpAdr[10]~0_combout\);

-- Location: FF_X80_Y8_N1
\R.curPC[10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[10]~0_combout\,
	asdata => \Add0~33_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(10));

-- Location: LABCELL_X81_Y6_N27
\Add0~37\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~37_sumout\ = SUM(( \R.curPC\(11) ) + ( GND ) + ( \Add0~34\ ))
-- \Add0~38\ = CARRY(( \R.curPC\(11) ) + ( GND ) + ( \Add0~34\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.curPC\(11),
	cin => \Add0~34\,
	sumout => \Add0~37_sumout\,
	cout => \Add0~38\);

-- Location: LABCELL_X83_Y6_N48
\R.regWriteData[11]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.regWriteData[11]~feeder_combout\ = ( \Add0~37_sumout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_Add0~37_sumout\,
	combout => \R.regWriteData[11]~feeder_combout\);

-- Location: LABCELL_X77_Y7_N45
\Selector21~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector21~0_combout\ = ( \Selector31~7_OTERM383\ & ( (!\R.aluData2\(3) & ((!\R.aluData2\(2) & (\ShiftRight1~32_OTERM21\)) # (\R.aluData2\(2) & ((\ShiftRight0~4_OTERM31\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000100010000010100010001000001010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(3),
	datab => \ALT_INV_ShiftRight1~32_OTERM21\,
	datac => \ALT_INV_ShiftRight0~4_OTERM31\,
	datad => \ALT_INV_R.aluData2\(2),
	dataf => \ALT_INV_Selector31~7_OTERM383\,
	combout => \Selector21~0_combout\);

-- Location: LABCELL_X71_Y6_N9
\Selector21~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector21~1_combout\ = ( !\R.aluData1\(11) & ( \R.aluOp.ALUOpOr~q\ & ( !\R.aluData2\(11) ) ) ) # ( \R.aluData1\(11) & ( !\R.aluOp.ALUOpOr~q\ & ( (!\R.aluData2\(11) & ((!\R.aluOp.ALUOpXor~DUPLICATE_q\))) # (\R.aluData2\(11) & 
-- (!\R.aluOp.ALUOpAnd~DUPLICATE_q\)) ) ) ) # ( !\R.aluData1\(11) & ( !\R.aluOp.ALUOpOr~q\ & ( (!\R.aluData2\(11)) # (!\R.aluOp.ALUOpXor~DUPLICATE_q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111110000111110100000101011110000111100000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpAnd~DUPLICATE_q\,
	datac => \ALT_INV_R.aluData2\(11),
	datad => \ALT_INV_R.aluOp.ALUOpXor~DUPLICATE_q\,
	datae => \ALT_INV_R.aluData1\(11),
	dataf => \ALT_INV_R.aluOp.ALUOpOr~q\,
	combout => \Selector21~1_combout\);

-- Location: FF_X71_Y7_N14
\ShiftRight0~7_NEW_REG232\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight0~7_RTM0235_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight0~7_OTERM233\);

-- Location: LABCELL_X71_Y6_N0
\Selector21~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector21~2_combout\ = ( \Selector31~6_OTERM381\ & ( \R.aluData1\(31) & ( (\Selector21~1_combout\ & (!\ShiftRight0~7_OTERM233\ & !\ShiftRight1~32_OTERM21\)) ) ) ) # ( !\Selector31~6_OTERM381\ & ( \R.aluData1\(31) & ( \Selector21~1_combout\ ) ) ) # ( 
-- \Selector31~6_OTERM381\ & ( !\R.aluData1\(31) & ( (\Selector21~1_combout\ & ((!\ShiftRight1~32_OTERM21\) # (\ShiftRight0~7_OTERM233\))) ) ) ) # ( !\Selector31~6_OTERM381\ & ( !\R.aluData1\(31) & ( \Selector21~1_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110011001100110000001100110011001100110011000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Selector21~1_combout\,
	datac => \ALT_INV_ShiftRight0~7_OTERM233\,
	datad => \ALT_INV_ShiftRight1~32_OTERM21\,
	datae => \ALT_INV_Selector31~6_OTERM381\,
	dataf => \ALT_INV_R.aluData1\(31),
	combout => \Selector21~2_combout\);

-- Location: LABCELL_X77_Y7_N36
\ShiftRight1~50\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~50_combout\ = ( \ShiftRight1~37_OTERM283\ & ( \ShiftRight1~30_OTERM39\ & ( (!\R.aluData2\(2) & (((\R.aluData2\(3)) # (\ShiftRight1~36_OTERM281\)))) # (\R.aluData2\(2) & (((!\R.aluData2\(3))) # (\ShiftRight1~31_OTERM45\))) ) ) ) # ( 
-- !\ShiftRight1~37_OTERM283\ & ( \ShiftRight1~30_OTERM39\ & ( (!\R.aluData2\(2) & (((\R.aluData2\(3)) # (\ShiftRight1~36_OTERM281\)))) # (\R.aluData2\(2) & (\ShiftRight1~31_OTERM45\ & ((\R.aluData2\(3))))) ) ) ) # ( \ShiftRight1~37_OTERM283\ & ( 
-- !\ShiftRight1~30_OTERM39\ & ( (!\R.aluData2\(2) & (((\ShiftRight1~36_OTERM281\ & !\R.aluData2\(3))))) # (\R.aluData2\(2) & (((!\R.aluData2\(3))) # (\ShiftRight1~31_OTERM45\))) ) ) ) # ( !\ShiftRight1~37_OTERM283\ & ( !\ShiftRight1~30_OTERM39\ & ( 
-- (!\R.aluData2\(2) & (((\ShiftRight1~36_OTERM281\ & !\R.aluData2\(3))))) # (\R.aluData2\(2) & (\ShiftRight1~31_OTERM45\ & ((\R.aluData2\(3))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000110000010001001111110001000100001100110111010011111111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~31_OTERM45\,
	datab => \ALT_INV_R.aluData2\(2),
	datac => \ALT_INV_ShiftRight1~36_OTERM281\,
	datad => \ALT_INV_R.aluData2\(3),
	datae => \ALT_INV_ShiftRight1~37_OTERM283\,
	dataf => \ALT_INV_ShiftRight1~30_OTERM39\,
	combout => \ShiftRight1~50_combout\);

-- Location: MLABCELL_X82_Y6_N18
\Selector21~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector21~3_combout\ = ( \Selector21~2_combout\ & ( \ShiftRight1~50_combout\ & ( (((\ShiftLeft0~15_combout\ & \Selector27~0_OTERM385\)) # (\Selector31~5_OTERM599\)) # (\Selector21~0_combout\) ) ) ) # ( !\Selector21~2_combout\ & ( 
-- \ShiftRight1~50_combout\ ) ) # ( \Selector21~2_combout\ & ( !\ShiftRight1~50_combout\ & ( ((\ShiftLeft0~15_combout\ & \Selector27~0_OTERM385\)) # (\Selector21~0_combout\) ) ) ) # ( !\Selector21~2_combout\ & ( !\ShiftRight1~50_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111001100110111011111111111111111110011111101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~15_combout\,
	datab => \ALT_INV_Selector21~0_combout\,
	datac => \ALT_INV_Selector31~5_OTERM599\,
	datad => \ALT_INV_Selector27~0_OTERM385\,
	datae => \ALT_INV_Selector21~2_combout\,
	dataf => \ALT_INV_ShiftRight1~50_combout\,
	combout => \Selector21~3_combout\);

-- Location: LABCELL_X83_Y6_N0
\Selector21~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector21~5_combout\ = ( \Add1~45_sumout\ & ( (((\Add2~45_sumout\ & \R.aluOp.ALUOpSub~q\)) # (\R.aluOp.ALUOpAdd~q\)) # (\Selector21~3_combout\) ) ) # ( !\Add1~45_sumout\ & ( ((\Add2~45_sumout\ & \R.aluOp.ALUOpSub~q\)) # (\Selector21~3_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001101110111001100110111011100111111011111110011111101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add2~45_sumout\,
	datab => \ALT_INV_Selector21~3_combout\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_R.aluOp.ALUOpSub~q\,
	dataf => \ALT_INV_Add1~45_sumout\,
	combout => \Selector21~5_combout\);

-- Location: FF_X83_Y6_N2
\R.aluRes[11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector21~5_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(11));

-- Location: LABCELL_X83_Y6_N51
\Comb:vRegWriteData[11]~1_RESYN1040\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[11]~1_RESYN1040_BDD1041\ = ( \Add2~45_sumout\ & ( ((!\R.aluCalc~q\ & (\R.aluRes\(11))) # (\R.aluCalc~q\ & ((\R.aluOp.ALUOpSub~q\)))) # (\R.memToReg~q\) ) ) # ( !\Add2~45_sumout\ & ( ((\R.aluRes\(11) & !\R.aluCalc~q\)) # 
-- (\R.memToReg~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101000011111111010100001111111101010011111111110101001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluRes\(11),
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_R.aluCalc~q\,
	datad => \ALT_INV_R.memToReg~q\,
	dataf => \ALT_INV_Add2~45_sumout\,
	combout => \Comb:vRegWriteData[11]~1_RESYN1040_BDD1041\);

-- Location: IOIBUF_X34_Y81_N92
\avm_d_readdata[19]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(19),
	o => \avm_d_readdata[19]~input_o\);

-- Location: LABCELL_X79_Y2_N54
\Comb:vRegWriteData[11]~1_RESYN1038\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[11]~1_RESYN1038_BDD1039\ = ( \avm_d_readdata[31]~input_o\ & ( \avm_d_readdata[19]~input_o\ & ( (!\R.memToReg~q\) # ((!\R.curInst\(12) & ((!\R.curInst\(14)))) # (\R.curInst\(12) & (!\R.curInst\(13)))) ) ) ) # ( 
-- !\avm_d_readdata[31]~input_o\ & ( \avm_d_readdata[19]~input_o\ & ( (!\R.memToReg~q\) # ((!\R.curInst\(13) & ((\R.curInst\(12)))) # (\R.curInst\(13) & (!\R.curInst\(14) & !\R.curInst\(12)))) ) ) ) # ( \avm_d_readdata[31]~input_o\ & ( 
-- !\avm_d_readdata[19]~input_o\ & ( (!\R.memToReg~q\) # ((!\R.curInst\(13) & (!\R.curInst\(14) & !\R.curInst\(12)))) ) ) ) # ( !\avm_d_readdata[31]~input_o\ & ( !\avm_d_readdata[19]~input_o\ & ( !\R.memToReg~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111100000000111111111000000011111111010010101111111111001010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(13),
	datab => \ALT_INV_R.curInst\(14),
	datac => \ALT_INV_R.curInst\(12),
	datad => \ALT_INV_R.memToReg~q\,
	datae => \ALT_INV_avm_d_readdata[31]~input_o\,
	dataf => \ALT_INV_avm_d_readdata[19]~input_o\,
	combout => \Comb:vRegWriteData[11]~1_RESYN1038_BDD1039\);

-- Location: LABCELL_X83_Y6_N42
\Comb:vRegWriteData[11]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[11]~1_combout\ = ( \Comb:vRegWriteData[11]~1_RESYN1040_BDD1041\ & ( \Comb:vRegWriteData[11]~1_RESYN1038_BDD1039\ ) ) # ( !\Comb:vRegWriteData[11]~1_RESYN1040_BDD1041\ & ( \Comb:vRegWriteData[11]~1_RESYN1038_BDD1039\ & ( (\R.aluCalc~q\ 
-- & (((\Add1~45_sumout\ & \R.aluOp.ALUOpAdd~q\)) # (\Selector21~3_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000001101111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add1~45_sumout\,
	datab => \ALT_INV_Selector21~3_combout\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_R.aluCalc~q\,
	datae => \ALT_INV_Comb:vRegWriteData[11]~1_RESYN1040_BDD1041\,
	dataf => \ALT_INV_Comb:vRegWriteData[11]~1_RESYN1038_BDD1039\,
	combout => \Comb:vRegWriteData[11]~1_combout\);

-- Location: FF_X83_Y6_N50
\R.regWriteData[11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \R.regWriteData[11]~feeder_combout\,
	asdata => \Comb:vRegWriteData[11]~1_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(11));

-- Location: FF_X66_Y2_N56
\RegFile[29][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(11),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][11]~q\);

-- Location: LABCELL_X73_Y2_N18
\Mux79~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux79~22_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[24][11]~q\))) # (\R.curInst\(15) & (\RegFile[25][11]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[26][11]~q\))) # (\R.curInst\(15) & (\RegFile[27][11]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[27][11]~q\,
	datab => \ALT_INV_RegFile[25][11]~q\,
	datac => \ALT_INV_RegFile[26][11]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][11]~q\,
	combout => \Mux79~22_combout\);

-- Location: LABCELL_X73_Y2_N54
\Mux79~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux79~9_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux79~22_combout\))))) # (\R.curInst\(17) & (((!\Mux79~22_combout\ & ((\RegFile[28][11]~q\))) # (\Mux79~22_combout\ & (\RegFile[29][11]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- (!\R.curInst\(17) & ((((\Mux79~22_combout\))))) # (\R.curInst\(17) & (((!\Mux79~22_combout\ & (\RegFile[30][11]~q\)) # (\Mux79~22_combout\ & ((\RegFile[31][11]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110111011101110111010101011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[29][11]~q\,
	datac => \ALT_INV_RegFile[30][11]~q\,
	datad => \ALT_INV_RegFile[31][11]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux79~22_combout\,
	datag => \ALT_INV_RegFile[28][11]~q\,
	combout => \Mux79~9_combout\);

-- Location: LABCELL_X61_Y2_N48
\Mux79~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux79~0_combout\ = ( \RegFile[7][11]~q\ & ( \R.curInst\(15) & ( (\RegFile[5][11]~q\) # (\R.curInst\(16)) ) ) ) # ( !\RegFile[7][11]~q\ & ( \R.curInst\(15) & ( (!\R.curInst\(16) & \RegFile[5][11]~q\) ) ) ) # ( \RegFile[7][11]~q\ & ( !\R.curInst\(15) & ( 
-- (!\R.curInst\(16) & (\RegFile[4][11]~q\)) # (\R.curInst\(16) & ((\RegFile[6][11]~q\))) ) ) ) # ( !\RegFile[7][11]~q\ & ( !\R.curInst\(15) & ( (!\R.curInst\(16) & (\RegFile[4][11]~q\)) # (\R.curInst\(16) & ((\RegFile[6][11]~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010011100100111001001110010011100000000101010100101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(16),
	datab => \ALT_INV_RegFile[4][11]~q\,
	datac => \ALT_INV_RegFile[6][11]~q\,
	datad => \ALT_INV_RegFile[5][11]~q\,
	datae => \ALT_INV_RegFile[7][11]~q\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux79~0_combout\);

-- Location: LABCELL_X61_Y2_N18
\Mux79~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux79~26_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (\RegFile[1][11]~q\ & (\R.curInst\(15)))) # (\R.curInst\(17) & (((\Mux79~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & ((!\R.curInst\(15) & (((\RegFile[2][11]~q\)))) # 
-- (\R.curInst\(15) & (\RegFile[3][11]~q\)))) # (\R.curInst\(17) & ((((\Mux79~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001100000011000100010000110011001111110011111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][11]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[2][11]~q\,
	datad => \ALT_INV_R.curInst\(15),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux79~0_combout\,
	datag => \ALT_INV_RegFile[1][11]~q\,
	combout => \Mux79~26_combout\);

-- Location: MLABCELL_X72_Y1_N18
\Mux79~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux79~18_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[16][11]~q\))) # (\R.curInst\(15) & (\RegFile[17][11]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[18][11]~q\))) # (\R.curInst\(15) & (\RegFile[19][11]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[17][11]~q\,
	datab => \ALT_INV_RegFile[19][11]~q\,
	datac => \ALT_INV_RegFile[18][11]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][11]~q\,
	combout => \Mux79~18_combout\);

-- Location: MLABCELL_X72_Y1_N12
\Mux79~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux79~5_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux79~18_combout\))))) # (\R.curInst\(17) & (((!\Mux79~18_combout\ & (\RegFile[20][11]~q\)) # (\Mux79~18_combout\ & ((\RegFile[21][11]~q\)))))) ) ) # ( \R.curInst\(16) & ( 
-- (!\R.curInst\(17) & ((((\Mux79~18_combout\))))) # (\R.curInst\(17) & (((!\Mux79~18_combout\ & ((\RegFile[22][11]~q\))) # (\Mux79~18_combout\ & (\RegFile[23][11]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110101010111111111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[23][11]~q\,
	datac => \ALT_INV_RegFile[22][11]~q\,
	datad => \ALT_INV_RegFile[21][11]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux79~18_combout\,
	datag => \ALT_INV_RegFile[20][11]~q\,
	combout => \Mux79~5_combout\);

-- Location: FF_X70_Y2_N44
\RegFile[11][11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[11][11]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][11]~q\);

-- Location: LABCELL_X70_Y2_N0
\Mux79~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux79~14_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[8][11]~q\))) # (\R.curInst\(15) & (\RegFile[9][11]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & (\RegFile[10][11]~q\)) # (\R.curInst\(15) & ((\RegFile[11][11]~q\))))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][11]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[10][11]~q\,
	datad => \ALT_INV_RegFile[11][11]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][11]~q\,
	combout => \Mux79~14_combout\);

-- Location: LABCELL_X73_Y2_N24
\Mux79~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux79~1_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux79~14_combout\)))) # (\R.curInst\(17) & ((!\Mux79~14_combout\ & ((\RegFile[12][11]~q\))) # (\Mux79~14_combout\ & (\RegFile[13][11]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux79~14_combout\)))) # (\R.curInst\(17) & ((!\Mux79~14_combout\ & ((\RegFile[14][11]~q\))) # (\Mux79~14_combout\ & (\RegFile[15][11]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][11]~q\,
	datab => \ALT_INV_RegFile[13][11]~q\,
	datac => \ALT_INV_RegFile[14][11]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux79~14_combout\,
	datag => \ALT_INV_RegFile[12][11]~q\,
	combout => \Mux79~1_combout\);

-- Location: LABCELL_X73_Y2_N15
\Mux79~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux79~13_combout\ = ( \Mux79~5_combout\ & ( \Mux79~1_combout\ & ( (!\R.curInst\(19) & (((\R.curInst\(18)) # (\Mux79~26_combout\)))) # (\R.curInst\(19) & (((!\R.curInst\(18))) # (\Mux79~9_combout\))) ) ) ) # ( !\Mux79~5_combout\ & ( \Mux79~1_combout\ & ( 
-- (!\R.curInst\(19) & (((\R.curInst\(18)) # (\Mux79~26_combout\)))) # (\R.curInst\(19) & (\Mux79~9_combout\ & ((\R.curInst\(18))))) ) ) ) # ( \Mux79~5_combout\ & ( !\Mux79~1_combout\ & ( (!\R.curInst\(19) & (((\Mux79~26_combout\ & !\R.curInst\(18))))) # 
-- (\R.curInst\(19) & (((!\R.curInst\(18))) # (\Mux79~9_combout\))) ) ) ) # ( !\Mux79~5_combout\ & ( !\Mux79~1_combout\ & ( (!\R.curInst\(19) & (((\Mux79~26_combout\ & !\R.curInst\(18))))) # (\R.curInst\(19) & (\Mux79~9_combout\ & ((\R.curInst\(18))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000110000010001001111110001000100001100110111010011111111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux79~9_combout\,
	datab => \ALT_INV_R.curInst\(19),
	datac => \ALT_INV_Mux79~26_combout\,
	datad => \ALT_INV_R.curInst\(18),
	datae => \ALT_INV_Mux79~5_combout\,
	dataf => \ALT_INV_Mux79~1_combout\,
	combout => \Mux79~13_combout\);

-- Location: LABCELL_X74_Y4_N57
\Mux243~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux243~0_combout\ = ( \Mux79~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC\(11)))) ) ) # ( !\Mux79~13_combout\ & ( (!\vAluSrc1~1_combout\ & (\vAluSrc1~2_combout\ & \R.curPC\(11))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000001010000000000000101010100000101010101010000010101010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluSrc1~1_combout\,
	datac => \ALT_INV_vAluSrc1~2_combout\,
	datad => \ALT_INV_R.curPC\(11),
	dataf => \ALT_INV_Mux79~13_combout\,
	combout => \Mux243~0_combout\);

-- Location: FF_X74_Y4_N29
\R.aluData1[11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux243~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData1\(11));

-- Location: LABCELL_X83_Y6_N12
\vAluRes~60\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~60_combout\ = ( !\R.aluCalc~q\ & ( (((\R.aluRes\(11)))) ) ) # ( \R.aluCalc~q\ & ( ((!\Add1~45_sumout\ & (\R.aluOp.ALUOpSub~q\ & ((\Add2~45_sumout\)))) # (\Add1~45_sumout\ & (((\R.aluOp.ALUOpSub~q\ & \Add2~45_sumout\)) # (\R.aluOp.ALUOpAdd~q\)))) 
-- # (\Selector21~3_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100001111000001011111111100001111000011110011011111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add1~45_sumout\,
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_Selector21~3_combout\,
	datae => \ALT_INV_R.aluCalc~q\,
	dataf => \ALT_INV_Add2~45_sumout\,
	datag => \ALT_INV_R.aluRes\(11),
	combout => \vAluRes~60_combout\);

-- Location: LABCELL_X80_Y4_N48
\Comb:vJumpAdr[11]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[11]~0_combout\ = ( \Add3~45_sumout\ & ( (!\Equal4~2_combout\) # (\vAluRes~60_combout\) ) ) # ( !\Add3~45_sumout\ & ( (\Equal4~2_combout\ & \vAluRes~60_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000110000001111001111110011111100111111001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Equal4~2_combout\,
	datac => \ALT_INV_vAluRes~60_combout\,
	dataf => \ALT_INV_Add3~45_sumout\,
	combout => \Comb:vJumpAdr[11]~0_combout\);

-- Location: FF_X80_Y4_N49
\R.curPC[11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[11]~0_combout\,
	asdata => \Add0~37_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(11));

-- Location: LABCELL_X81_Y6_N30
\Add0~41\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~41_sumout\ = SUM(( \R.curPC\(12) ) + ( GND ) + ( \Add0~38\ ))
-- \Add0~42\ = CARRY(( \R.curPC\(12) ) + ( GND ) + ( \Add0~38\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.curPC\(12),
	cin => \Add0~38\,
	sumout => \Add0~41_sumout\,
	cout => \Add0~42\);

-- Location: LABCELL_X81_Y4_N12
\R.regWriteData[12]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.regWriteData[12]~feeder_combout\ = ( \Add0~41_sumout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_Add0~41_sumout\,
	combout => \R.regWriteData[12]~feeder_combout\);

-- Location: LABCELL_X81_Y4_N15
\Comb:vRegWriteData[12]~1_RESYN1088\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[12]~1_RESYN1088_BDD1089\ = ( \R.aluCalc~q\ & ( ((\R.aluOp.ALUOpSub~q\ & \Add2~49_sumout\)) # (\R.memToReg~q\) ) ) # ( !\R.aluCalc~q\ & ( (\R.aluRes\(12)) # (\R.memToReg~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001111111111001100111111111100110111001101110011011100110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datab => \ALT_INV_R.memToReg~q\,
	datac => \ALT_INV_Add2~49_sumout\,
	datad => \ALT_INV_R.aluRes\(12),
	dataf => \ALT_INV_R.aluCalc~q\,
	combout => \Comb:vRegWriteData[12]~1_RESYN1088_BDD1089\);

-- Location: IOIBUF_X62_Y0_N18
\avm_d_readdata[20]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(20),
	o => \avm_d_readdata[20]~input_o\);

-- Location: LABCELL_X79_Y2_N51
\Comb:vRegWriteData[12]~1_RESYN1086\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[12]~1_RESYN1086_BDD1087\ = ( \avm_d_readdata[31]~input_o\ & ( \avm_d_readdata[20]~input_o\ & ( (!\R.memToReg~q\) # ((!\R.curInst\(12) & ((!\R.curInst\(14)))) # (\R.curInst\(12) & (!\R.curInst\(13)))) ) ) ) # ( 
-- !\avm_d_readdata[31]~input_o\ & ( \avm_d_readdata[20]~input_o\ & ( (!\R.memToReg~q\) # ((!\R.curInst\(13) & ((\R.curInst\(12)))) # (\R.curInst\(13) & (!\R.curInst\(14) & !\R.curInst\(12)))) ) ) ) # ( \avm_d_readdata[31]~input_o\ & ( 
-- !\avm_d_readdata[20]~input_o\ & ( (!\R.memToReg~q\) # ((!\R.curInst\(13) & (!\R.curInst\(14) & !\R.curInst\(12)))) ) ) ) # ( !\avm_d_readdata[31]~input_o\ & ( !\avm_d_readdata[20]~input_o\ & ( !\R.memToReg~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111000011110000111110001111000011110100111110101111110011111010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(13),
	datab => \ALT_INV_R.curInst\(14),
	datac => \ALT_INV_R.memToReg~q\,
	datad => \ALT_INV_R.curInst\(12),
	datae => \ALT_INV_avm_d_readdata[31]~input_o\,
	dataf => \ALT_INV_avm_d_readdata[20]~input_o\,
	combout => \Comb:vRegWriteData[12]~1_RESYN1086_BDD1087\);

-- Location: LABCELL_X81_Y4_N54
\Comb:vRegWriteData[12]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[12]~1_combout\ = ( \Comb:vRegWriteData[12]~1_RESYN1086_BDD1087\ & ( \Selector20~3_combout\ & ( ((\R.aluCalc~q\ & (\Add1~49_sumout\ & \R.aluOp.ALUOpAdd~q\))) # (\Comb:vRegWriteData[12]~1_RESYN1088_BDD1089\) ) ) ) # ( 
-- \Comb:vRegWriteData[12]~1_RESYN1086_BDD1087\ & ( !\Selector20~3_combout\ & ( (\Comb:vRegWriteData[12]~1_RESYN1088_BDD1089\) # (\R.aluCalc~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010101011111111100000000000000000000000111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluCalc~q\,
	datab => \ALT_INV_Add1~49_sumout\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_Comb:vRegWriteData[12]~1_RESYN1088_BDD1089\,
	datae => \ALT_INV_Comb:vRegWriteData[12]~1_RESYN1086_BDD1087\,
	dataf => \ALT_INV_Selector20~3_combout\,
	combout => \Comb:vRegWriteData[12]~1_combout\);

-- Location: FF_X81_Y4_N14
\R.regWriteData[12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \R.regWriteData[12]~feeder_combout\,
	asdata => \Comb:vRegWriteData[12]~1_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(12));

-- Location: LABCELL_X68_Y8_N30
\RegFile[13][12]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[13][12]~feeder_combout\ = ( \R.regWriteData\(12) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(12),
	combout => \RegFile[13][12]~feeder_combout\);

-- Location: FF_X68_Y8_N31
\RegFile[13][12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[13][12]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][12]~q\);

-- Location: LABCELL_X66_Y8_N6
\Mux78~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux78~14_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[8][12]~q\))) # (\R.curInst\(15) & (\RegFile[9][12]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & (\RegFile[10][12]~q\)) # (\R.curInst\(15) & ((\RegFile[11][12]~q\))))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][12]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[10][12]~q\,
	datad => \ALT_INV_RegFile[11][12]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][12]~q\,
	combout => \Mux78~14_combout\);

-- Location: LABCELL_X66_Y8_N42
\Mux78~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux78~1_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux78~14_combout\)))) # (\R.curInst\(17) & ((!\Mux78~14_combout\ & ((\RegFile[12][12]~q\))) # (\Mux78~14_combout\ & (\RegFile[13][12]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux78~14_combout\)))) # (\R.curInst\(17) & ((!\Mux78~14_combout\ & ((\RegFile[14][12]~q\))) # (\Mux78~14_combout\ & (\RegFile[15][12]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][12]~q\,
	datab => \ALT_INV_RegFile[15][12]~q\,
	datac => \ALT_INV_RegFile[14][12]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux78~14_combout\,
	datag => \ALT_INV_RegFile[12][12]~q\,
	combout => \Mux78~1_combout\);

-- Location: MLABCELL_X65_Y6_N0
\Mux78~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux78~0_combout\ = ( \RegFile[7][12]~q\ & ( \R.curInst\(15) & ( (\R.curInst\(16)) # (\RegFile[5][12]~q\) ) ) ) # ( !\RegFile[7][12]~q\ & ( \R.curInst\(15) & ( (\RegFile[5][12]~q\ & !\R.curInst\(16)) ) ) ) # ( \RegFile[7][12]~q\ & ( !\R.curInst\(15) & ( 
-- (!\R.curInst\(16) & ((\RegFile[4][12]~q\))) # (\R.curInst\(16) & (\RegFile[6][12]~q\)) ) ) ) # ( !\RegFile[7][12]~q\ & ( !\R.curInst\(15) & ( (!\R.curInst\(16) & ((\RegFile[4][12]~q\))) # (\R.curInst\(16) & (\RegFile[6][12]~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001111110011000000111111001101010000010100000101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[5][12]~q\,
	datab => \ALT_INV_RegFile[6][12]~q\,
	datac => \ALT_INV_R.curInst\(16),
	datad => \ALT_INV_RegFile[4][12]~q\,
	datae => \ALT_INV_RegFile[7][12]~q\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux78~0_combout\);

-- Location: FF_X65_Y6_N55
\RegFile[2][12]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(12),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][12]~DUPLICATE_q\);

-- Location: LABCELL_X70_Y8_N33
\Mux78~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux78~26_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((\RegFile[1][12]~q\ & ((\R.curInst\(15))))))) # (\R.curInst\(17) & (\Mux78~0_combout\)) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & (\RegFile[2][12]~DUPLICATE_q\)) 
-- # (\R.curInst\(15) & ((\RegFile[3][12]~q\)))))) # (\R.curInst\(17) & (\Mux78~0_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0001000100010001000110110001101100011011000110110001000110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_Mux78~0_combout\,
	datac => \ALT_INV_RegFile[2][12]~DUPLICATE_q\,
	datad => \ALT_INV_RegFile[3][12]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[1][12]~q\,
	combout => \Mux78~26_combout\);

-- Location: LABCELL_X68_Y8_N36
\Mux78~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux78~18_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[16][12]~q\))) # (\R.curInst\(15) & (\RegFile[17][12]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[18][12]~q\))) # (\R.curInst\(15) & (\RegFile[19][12]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[19][12]~q\,
	datab => \ALT_INV_RegFile[17][12]~q\,
	datac => \ALT_INV_RegFile[18][12]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][12]~q\,
	combout => \Mux78~18_combout\);

-- Location: LABCELL_X70_Y8_N36
\Mux78~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux78~5_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux78~18_combout\))))) # (\R.curInst\(17) & (((!\Mux78~18_combout\ & (\RegFile[20][12]~q\)) # (\Mux78~18_combout\ & ((\RegFile[21][12]~q\)))))) ) ) # ( \R.curInst\(16) & ( 
-- (!\R.curInst\(17) & ((((\Mux78~18_combout\))))) # (\R.curInst\(17) & (((!\Mux78~18_combout\ & ((\RegFile[22][12]~q\))) # (\Mux78~18_combout\ & (\RegFile[23][12]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110101010111111111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[23][12]~q\,
	datac => \ALT_INV_RegFile[22][12]~q\,
	datad => \ALT_INV_RegFile[21][12]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux78~18_combout\,
	datag => \ALT_INV_RegFile[20][12]~q\,
	combout => \Mux78~5_combout\);

-- Location: MLABCELL_X65_Y4_N48
\Mux78~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux78~22_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[24][12]~q\))) # (\R.curInst\(15) & (\RegFile[25][12]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & (\RegFile[26][12]~q\)) # (\R.curInst\(15) & ((\RegFile[27][12]~q\))))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[25][12]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[26][12]~q\,
	datad => \ALT_INV_RegFile[27][12]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][12]~q\,
	combout => \Mux78~22_combout\);

-- Location: MLABCELL_X65_Y4_N0
\Mux78~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux78~9_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux78~22_combout\)))) # (\R.curInst\(17) & ((!\Mux78~22_combout\ & (\RegFile[28][12]~q\)) # (\Mux78~22_combout\ & ((\RegFile[29][12]~q\)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) 
-- & ((((\Mux78~22_combout\))))) # (\R.curInst\(17) & (((!\Mux78~22_combout\ & ((\RegFile[30][12]~q\))) # (\Mux78~22_combout\ & (\RegFile[31][12]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111001100111111111101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][12]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[30][12]~q\,
	datad => \ALT_INV_RegFile[29][12]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux78~22_combout\,
	datag => \ALT_INV_RegFile[28][12]~q\,
	combout => \Mux78~9_combout\);

-- Location: LABCELL_X70_Y8_N48
\Mux78~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux78~13_combout\ = ( \Mux78~5_combout\ & ( \Mux78~9_combout\ & ( ((!\R.curInst\(18) & ((\Mux78~26_combout\))) # (\R.curInst\(18) & (\Mux78~1_combout\))) # (\R.curInst\(19)) ) ) ) # ( !\Mux78~5_combout\ & ( \Mux78~9_combout\ & ( (!\R.curInst\(19) & 
-- ((!\R.curInst\(18) & ((\Mux78~26_combout\))) # (\R.curInst\(18) & (\Mux78~1_combout\)))) # (\R.curInst\(19) & (((\R.curInst\(18))))) ) ) ) # ( \Mux78~5_combout\ & ( !\Mux78~9_combout\ & ( (!\R.curInst\(19) & ((!\R.curInst\(18) & ((\Mux78~26_combout\))) # 
-- (\R.curInst\(18) & (\Mux78~1_combout\)))) # (\R.curInst\(19) & (((!\R.curInst\(18))))) ) ) ) # ( !\Mux78~5_combout\ & ( !\Mux78~9_combout\ & ( (!\R.curInst\(19) & ((!\R.curInst\(18) & ((\Mux78~26_combout\))) # (\R.curInst\(18) & (\Mux78~1_combout\)))) ) ) 
-- )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101000100010010111110010001000001010011101110101111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(19),
	datab => \ALT_INV_Mux78~1_combout\,
	datac => \ALT_INV_Mux78~26_combout\,
	datad => \ALT_INV_R.curInst\(18),
	datae => \ALT_INV_Mux78~5_combout\,
	dataf => \ALT_INV_Mux78~9_combout\,
	combout => \Mux78~13_combout\);

-- Location: LABCELL_X70_Y8_N18
\Mux242~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux242~0_combout\ = ( !\vAluSrc1~1_combout\ & ( \Mux78~13_combout\ & ( (!\vAluSrc1~2_combout\) # (\R.curPC\(12)) ) ) ) # ( !\vAluSrc1~1_combout\ & ( !\Mux78~13_combout\ & ( (\R.curPC\(12) & \vAluSrc1~2_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010101000000000000000011111111010101010000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curPC\(12),
	datad => \ALT_INV_vAluSrc1~2_combout\,
	datae => \ALT_INV_vAluSrc1~1_combout\,
	dataf => \ALT_INV_Mux78~13_combout\,
	combout => \Mux242~0_combout\);

-- Location: FF_X74_Y6_N22
\R.aluData1[12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \Mux242~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData1\(12));

-- Location: LABCELL_X81_Y4_N39
\Selector20~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector20~4_combout\ = ( \Add1~49_sumout\ & ( ((\R.aluOp.ALUOpSub~q\ & \Add2~49_sumout\)) # (\R.aluOp.ALUOpAdd~q\) ) ) # ( !\Add1~49_sumout\ & ( (\R.aluOp.ALUOpSub~q\ & \Add2~49_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011010101110101011100000011000000110101011101010111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_Add2~49_sumout\,
	datae => \ALT_INV_Add1~49_sumout\,
	combout => \Selector20~4_combout\);

-- Location: LABCELL_X81_Y4_N24
\Comb:vJumpAdr[12]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[12]~0_combout\ = ( \Equal4~2_combout\ & ( \Add3~49_sumout\ & ( (!\R.aluCalc~q\ & (((\R.aluRes\(12))))) # (\R.aluCalc~q\ & (((!\Selector20~3_combout\)) # (\Selector20~4_combout\))) ) ) ) # ( !\Equal4~2_combout\ & ( \Add3~49_sumout\ ) ) # ( 
-- \Equal4~2_combout\ & ( !\Add3~49_sumout\ & ( (!\R.aluCalc~q\ & (((\R.aluRes\(12))))) # (\R.aluCalc~q\ & (((!\Selector20~3_combout\)) # (\Selector20~4_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010100011111101111111111111111110101000111111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluCalc~q\,
	datab => \ALT_INV_Selector20~4_combout\,
	datac => \ALT_INV_Selector20~3_combout\,
	datad => \ALT_INV_R.aluRes\(12),
	datae => \ALT_INV_Equal4~2_combout\,
	dataf => \ALT_INV_Add3~49_sumout\,
	combout => \Comb:vJumpAdr[12]~0_combout\);

-- Location: FF_X81_Y4_N25
\R.curPC[12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[12]~0_combout\,
	asdata => \Add0~41_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(12));

-- Location: MLABCELL_X78_Y8_N15
\R.regWriteData[13]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.regWriteData[13]~feeder_combout\ = \Add0~45_sumout\

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Add0~45_sumout\,
	combout => \R.regWriteData[13]~feeder_combout\);

-- Location: FF_X71_Y6_N17
\R.aluData2[13]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \NxR.aluData2[13]~10_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData2[13]~DUPLICATE_q\);

-- Location: LABCELL_X71_Y6_N30
\Selector19~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector19~2_combout\ = ( !\R.aluData1\(13) & ( \R.aluOp.ALUOpOr~q\ & ( !\R.aluData2[13]~DUPLICATE_q\ ) ) ) # ( \R.aluData1\(13) & ( !\R.aluOp.ALUOpOr~q\ & ( (!\R.aluData2[13]~DUPLICATE_q\ & (!\R.aluOp.ALUOpXor~DUPLICATE_q\)) # 
-- (\R.aluData2[13]~DUPLICATE_q\ & ((!\R.aluOp.ALUOpAnd~DUPLICATE_q\))) ) ) ) # ( !\R.aluData1\(13) & ( !\R.aluOp.ALUOpOr~q\ & ( (!\R.aluOp.ALUOpXor~DUPLICATE_q\) # (!\R.aluData2[13]~DUPLICATE_q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1110111011101110101110001011100011001100110011000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpXor~DUPLICATE_q\,
	datab => \ALT_INV_R.aluData2[13]~DUPLICATE_q\,
	datac => \ALT_INV_R.aluOp.ALUOpAnd~DUPLICATE_q\,
	datae => \ALT_INV_R.aluData1\(13),
	dataf => \ALT_INV_R.aluOp.ALUOpOr~q\,
	combout => \Selector19~2_combout\);

-- Location: MLABCELL_X78_Y9_N0
\ShiftRight1~52\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~52_combout\ = ( \ShiftRight1~11_OTERM35\ & ( \R.aluData2\(3) & ( (!\R.aluData2\(2)) # (\ShiftRight1~12_OTERM57\) ) ) ) # ( !\ShiftRight1~11_OTERM35\ & ( \R.aluData2\(3) & ( (\ShiftRight1~12_OTERM57\ & \R.aluData2\(2)) ) ) ) # ( 
-- \ShiftRight1~11_OTERM35\ & ( !\R.aluData2\(3) & ( (!\R.aluData2\(2) & ((\ShiftRight1~18_OTERM269\))) # (\R.aluData2\(2) & (\ShiftRight1~10_OTERM265\)) ) ) ) # ( !\ShiftRight1~11_OTERM35\ & ( !\R.aluData2\(3) & ( (!\R.aluData2\(2) & 
-- ((\ShiftRight1~18_OTERM269\))) # (\R.aluData2\(2) & (\ShiftRight1~10_OTERM265\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111101010101000011110101010100000000001100111111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~10_OTERM265\,
	datab => \ALT_INV_ShiftRight1~12_OTERM57\,
	datac => \ALT_INV_ShiftRight1~18_OTERM269\,
	datad => \ALT_INV_R.aluData2\(2),
	datae => \ALT_INV_ShiftRight1~11_OTERM35\,
	dataf => \ALT_INV_R.aluData2\(3),
	combout => \ShiftRight1~52_combout\);

-- Location: LABCELL_X74_Y5_N24
\Selector19~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector19~0_combout\ = ( !\NxR.aluData2[1]~17_combout\ & ( \NxR.aluData2[0]~16_combout\ & ( (\Mux224~0_combout\ & \R.aluOp.ALUOpSRL_OTERM361\) ) ) ) # ( \NxR.aluData2[1]~17_combout\ & ( !\NxR.aluData2[0]~16_combout\ & ( (\Mux223~0_combout\ & 
-- \R.aluOp.ALUOpSRL_OTERM361\) ) ) ) # ( !\NxR.aluData2[1]~17_combout\ & ( !\NxR.aluData2[0]~16_combout\ & ( (\R.aluOp.ALUOpSRL_OTERM361\ & \Mux225~0_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000001111000000110000001100000101000001010000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux224~0_combout\,
	datab => \ALT_INV_Mux223~0_combout\,
	datac => \ALT_INV_R.aluOp.ALUOpSRL_OTERM361\,
	datad => \ALT_INV_Mux225~0_combout\,
	datae => \ALT_INV_NxR.aluData2[1]~17_combout\,
	dataf => \ALT_INV_NxR.aluData2[0]~16_combout\,
	combout => \Selector19~0_combout\);

-- Location: FF_X74_Y5_N25
\Selector19~1_OTERM751_NEW_REG802\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector19~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector19~1_OTERM751_OTERM803\);

-- Location: LABCELL_X79_Y7_N12
\Selector19~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector19~1_combout\ = ( \R.aluOp.ALUOpSRA~q\ & ( \R.aluData2\(4) & ( (!\ShiftRight0~7_OTERM233DUPLICATE_q\ & (((\ShiftRight1~13_OTERM15\)) # (\Selector19~1_OTERM751_OTERM803\))) # (\ShiftRight0~7_OTERM233DUPLICATE_q\ & (((\R.aluData1\(31))))) ) ) ) # ( 
-- !\R.aluOp.ALUOpSRA~q\ & ( \R.aluData2\(4) & ( (\Selector19~1_OTERM751_OTERM803\ & !\ShiftRight0~7_OTERM233DUPLICATE_q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000001010101000000000101111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector19~1_OTERM751_OTERM803\,
	datab => \ALT_INV_R.aluData1\(31),
	datac => \ALT_INV_ShiftRight1~13_OTERM15\,
	datad => \ALT_INV_ShiftRight0~7_OTERM233DUPLICATE_q\,
	datae => \ALT_INV_R.aluOp.ALUOpSRA~q\,
	dataf => \ALT_INV_R.aluData2\(4),
	combout => \Selector19~1_combout\);

-- Location: LABCELL_X79_Y7_N54
\Selector19~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector19~3_combout\ = ( \Selector31~5_OTERM599\ & ( \Selector19~1_combout\ ) ) # ( !\Selector31~5_OTERM599\ & ( \Selector19~1_combout\ ) ) # ( \Selector31~5_OTERM599\ & ( !\Selector19~1_combout\ & ( (!\Selector19~2_combout\) # 
-- (((\ShiftLeft0~19_combout\ & \Selector27~0_OTERM385\)) # (\ShiftRight1~52_combout\)) ) ) ) # ( !\Selector31~5_OTERM599\ & ( !\Selector19~1_combout\ & ( (!\Selector19~2_combout\) # ((\ShiftLeft0~19_combout\ & \Selector27~0_OTERM385\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1100110111001101110011011111111111111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~19_combout\,
	datab => \ALT_INV_Selector19~2_combout\,
	datac => \ALT_INV_Selector27~0_OTERM385\,
	datad => \ALT_INV_ShiftRight1~52_combout\,
	datae => \ALT_INV_Selector31~5_OTERM599\,
	dataf => \ALT_INV_Selector19~1_combout\,
	combout => \Selector19~3_combout\);

-- Location: MLABCELL_X78_Y8_N6
\Selector19~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector19~5_combout\ = ( \Selector19~3_combout\ & ( \R.aluOp.ALUOpAdd~q\ ) ) # ( !\Selector19~3_combout\ & ( \R.aluOp.ALUOpAdd~q\ & ( ((\R.aluOp.ALUOpSub~q\ & \Add2~53_sumout\)) # (\Add1~53_sumout\) ) ) ) # ( \Selector19~3_combout\ & ( 
-- !\R.aluOp.ALUOpAdd~q\ ) ) # ( !\Selector19~3_combout\ & ( !\R.aluOp.ALUOpAdd~q\ & ( (\R.aluOp.ALUOpSub~q\ & \Add2~53_sumout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100010001111111111111111100010001111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datab => \ALT_INV_Add2~53_sumout\,
	datad => \ALT_INV_Add1~53_sumout\,
	datae => \ALT_INV_Selector19~3_combout\,
	dataf => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	combout => \Selector19~5_combout\);

-- Location: FF_X78_Y8_N7
\R.aluRes[13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector19~5_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(13));

-- Location: LABCELL_X79_Y8_N33
\Comb:vRegWriteData[13]~1_RESYN1044\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[13]~1_RESYN1044_BDD1045\ = ( \R.memToReg~q\ & ( \Add2~53_sumout\ ) ) # ( !\R.memToReg~q\ & ( \Add2~53_sumout\ & ( (!\R.aluCalc~q\ & (\R.aluRes\(13))) # (\R.aluCalc~q\ & ((\R.aluOp.ALUOpSub~q\))) ) ) ) # ( \R.memToReg~q\ & ( 
-- !\Add2~53_sumout\ ) ) # ( !\R.memToReg~q\ & ( !\Add2~53_sumout\ & ( (\R.aluRes\(13) & !\R.aluCalc~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101000001010000111111111111111101010000010111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluRes\(13),
	datac => \ALT_INV_R.aluCalc~q\,
	datad => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datae => \ALT_INV_R.memToReg~q\,
	dataf => \ALT_INV_Add2~53_sumout\,
	combout => \Comb:vRegWriteData[13]~1_RESYN1044_BDD1045\);

-- Location: IOIBUF_X36_Y0_N18
\avm_d_readdata[21]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(21),
	o => \avm_d_readdata[21]~input_o\);

-- Location: LABCELL_X79_Y2_N57
\Comb:vRegWriteData[13]~1_RESYN1042\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[13]~1_RESYN1042_BDD1043\ = ( \avm_d_readdata[31]~input_o\ & ( \avm_d_readdata[21]~input_o\ & ( (!\R.memToReg~q\) # ((!\R.curInst\(12) & ((!\R.curInst\(14)))) # (\R.curInst\(12) & (!\R.curInst\(13)))) ) ) ) # ( 
-- !\avm_d_readdata[31]~input_o\ & ( \avm_d_readdata[21]~input_o\ & ( (!\R.memToReg~q\) # ((!\R.curInst\(13) & ((\R.curInst\(12)))) # (\R.curInst\(13) & (!\R.curInst\(14) & !\R.curInst\(12)))) ) ) ) # ( \avm_d_readdata[31]~input_o\ & ( 
-- !\avm_d_readdata[21]~input_o\ & ( (!\R.memToReg~q\) # ((!\R.curInst\(13) & (!\R.curInst\(14) & !\R.curInst\(12)))) ) ) ) # ( !\avm_d_readdata[31]~input_o\ & ( !\avm_d_readdata[21]~input_o\ & ( !\R.memToReg~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111000011110000111110001111000011110100111110101111110011111010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(13),
	datab => \ALT_INV_R.curInst\(14),
	datac => \ALT_INV_R.memToReg~q\,
	datad => \ALT_INV_R.curInst\(12),
	datae => \ALT_INV_avm_d_readdata[31]~input_o\,
	dataf => \ALT_INV_avm_d_readdata[21]~input_o\,
	combout => \Comb:vRegWriteData[13]~1_RESYN1042_BDD1043\);

-- Location: MLABCELL_X78_Y8_N36
\Comb:vRegWriteData[13]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[13]~1_combout\ = ( \Selector19~3_combout\ & ( \Comb:vRegWriteData[13]~1_RESYN1042_BDD1043\ & ( (\Comb:vRegWriteData[13]~1_RESYN1044_BDD1045\) # (\R.aluCalc~q\) ) ) ) # ( !\Selector19~3_combout\ & ( 
-- \Comb:vRegWriteData[13]~1_RESYN1042_BDD1043\ & ( ((\R.aluCalc~q\ & (\R.aluOp.ALUOpAdd~q\ & \Add1~53_sumout\))) # (\Comb:vRegWriteData[13]~1_RESYN1044_BDD1045\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000001111000111110101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluCalc~q\,
	datab => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datac => \ALT_INV_Comb:vRegWriteData[13]~1_RESYN1044_BDD1045\,
	datad => \ALT_INV_Add1~53_sumout\,
	datae => \ALT_INV_Selector19~3_combout\,
	dataf => \ALT_INV_Comb:vRegWriteData[13]~1_RESYN1042_BDD1043\,
	combout => \Comb:vRegWriteData[13]~1_combout\);

-- Location: FF_X78_Y8_N17
\R.regWriteData[13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \R.regWriteData[13]~feeder_combout\,
	asdata => \Comb:vRegWriteData[13]~1_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(13));

-- Location: LABCELL_X71_Y2_N54
\RegFile[29][13]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[29][13]~feeder_combout\ = ( \R.regWriteData\(13) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(13),
	combout => \RegFile[29][13]~feeder_combout\);

-- Location: FF_X71_Y2_N55
\RegFile[29][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[29][13]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][13]~q\);

-- Location: FF_X73_Y2_N20
\RegFile[30][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(13),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][13]~q\);

-- Location: FF_X73_Y2_N38
\RegFile[31][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(13),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][13]~q\);

-- Location: FF_X67_Y2_N20
\RegFile[27][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(13),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][13]~q\);

-- Location: FF_X67_Y2_N8
\RegFile[25][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(13),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][13]~q\);

-- Location: FF_X67_Y2_N50
\RegFile[26][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(13),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][13]~q\);

-- Location: FF_X59_Y2_N44
\RegFile[24][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(13),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][13]~q\);

-- Location: LABCELL_X67_Y2_N6
\Mux109~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux109~22_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[24][13]~q\))) # (\R.curInst\(20) & (\RegFile[25][13]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[26][13]~q\))) # (\R.curInst\(20) & (\RegFile[27][13]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[27][13]~q\,
	datab => \ALT_INV_RegFile[25][13]~q\,
	datac => \ALT_INV_RegFile[26][13]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][13]~q\,
	combout => \Mux109~22_combout\);

-- Location: LABCELL_X73_Y2_N33
\RegFile[28][13]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[28][13]~feeder_combout\ = ( \R.regWriteData\(13) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(13),
	combout => \RegFile[28][13]~feeder_combout\);

-- Location: FF_X73_Y2_N34
\RegFile[28][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[28][13]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][13]~q\);

-- Location: LABCELL_X71_Y2_N21
\Mux109~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux109~9_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux109~22_combout\))))) # (\R.curInst\(22) & (((!\Mux109~22_combout\ & ((\RegFile[28][13]~q\))) # (\Mux109~22_combout\ & (\RegFile[29][13]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- (!\R.curInst\(22) & ((((\Mux109~22_combout\))))) # (\R.curInst\(22) & (((!\Mux109~22_combout\ & (\RegFile[30][13]~q\)) # (\Mux109~22_combout\ & ((\RegFile[31][13]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110111011101110111010101011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[29][13]~q\,
	datac => \ALT_INV_RegFile[30][13]~q\,
	datad => \ALT_INV_RegFile[31][13]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux109~22_combout\,
	datag => \ALT_INV_RegFile[28][13]~q\,
	combout => \Mux109~9_combout\);

-- Location: FF_X71_Y2_N44
\RegFile[13][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(13),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][13]~q\);

-- Location: FF_X62_Y2_N23
\RegFile[14][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(13),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][13]~q\);

-- Location: FF_X70_Y2_N26
\RegFile[15][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(13),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][13]~q\);

-- Location: FF_X70_Y2_N20
\RegFile[11][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(13),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][13]~q\);

-- Location: LABCELL_X73_Y1_N18
\RegFile[10][13]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[10][13]~feeder_combout\ = ( \R.regWriteData\(13) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(13),
	combout => \RegFile[10][13]~feeder_combout\);

-- Location: FF_X73_Y1_N19
\RegFile[10][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[10][13]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][13]~q\);

-- Location: FF_X70_Y2_N38
\RegFile[9][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(13),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][13]~q\);

-- Location: FF_X68_Y5_N31
\RegFile[8][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(13),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][13]~q\);

-- Location: LABCELL_X70_Y2_N36
\Mux109~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux109~14_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & (\RegFile[8][13]~q\)) # (\R.curInst\(20) & ((\RegFile[9][13]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & ((\RegFile[10][13]~q\))) # (\R.curInst\(20) & (\RegFile[11][13]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110000110011111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[11][13]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[10][13]~q\,
	datad => \ALT_INV_RegFile[9][13]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][13]~q\,
	combout => \Mux109~14_combout\);

-- Location: LABCELL_X62_Y2_N42
\RegFile[12][13]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[12][13]~feeder_combout\ = \R.regWriteData\(13)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.regWriteData\(13),
	combout => \RegFile[12][13]~feeder_combout\);

-- Location: FF_X62_Y2_N44
\RegFile[12][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[12][13]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][13]~q\);

-- Location: LABCELL_X71_Y2_N42
\Mux109~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux109~1_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux109~14_combout\))))) # (\R.curInst\(22) & (((!\Mux109~14_combout\ & ((\RegFile[12][13]~q\))) # (\Mux109~14_combout\ & (\RegFile[13][13]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux109~14_combout\)))) # (\R.curInst\(22) & ((!\Mux109~14_combout\ & (\RegFile[14][13]~q\)) # (\Mux109~14_combout\ & ((\RegFile[15][13]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][13]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[14][13]~q\,
	datad => \ALT_INV_RegFile[15][13]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux109~14_combout\,
	datag => \ALT_INV_RegFile[12][13]~q\,
	combout => \Mux109~1_combout\);

-- Location: FF_X73_Y3_N8
\RegFile[3][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(13),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][13]~q\);

-- Location: FF_X72_Y3_N20
\RegFile[2][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(13),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][13]~q\);

-- Location: FF_X67_Y5_N55
\RegFile[4][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(13),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][13]~q\);

-- Location: FF_X73_Y3_N44
\RegFile[7][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(13),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][13]~q\);

-- Location: FF_X73_Y3_N29
\RegFile[6][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(13),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][13]~q\);

-- Location: FF_X72_Y3_N13
\RegFile[5][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(13),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][13]~q\);

-- Location: MLABCELL_X72_Y3_N12
\Mux109~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux109~0_combout\ = ( \RegFile[5][13]~q\ & ( \R.curInst\(20) & ( (!\R.curInst\(21)) # (\RegFile[7][13]~q\) ) ) ) # ( !\RegFile[5][13]~q\ & ( \R.curInst\(20) & ( (\RegFile[7][13]~q\ & \R.curInst\(21)) ) ) ) # ( \RegFile[5][13]~q\ & ( !\R.curInst\(20) & ( 
-- (!\R.curInst\(21) & (\RegFile[4][13]~q\)) # (\R.curInst\(21) & ((\RegFile[6][13]~q\))) ) ) ) # ( !\RegFile[5][13]~q\ & ( !\R.curInst\(20) & ( (!\R.curInst\(21) & (\RegFile[4][13]~q\)) # (\R.curInst\(21) & ((\RegFile[6][13]~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101000001011111010100000101111100000011000000111111001111110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[4][13]~q\,
	datab => \ALT_INV_RegFile[7][13]~q\,
	datac => \ALT_INV_R.curInst\(21),
	datad => \ALT_INV_RegFile[6][13]~q\,
	datae => \ALT_INV_RegFile[5][13]~q\,
	dataf => \ALT_INV_R.curInst\(20),
	combout => \Mux109~0_combout\);

-- Location: FF_X72_Y3_N31
\RegFile[1][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(13),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][13]~q\);

-- Location: MLABCELL_X72_Y3_N18
\Mux109~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux109~26_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((\RegFile[1][13]~q\ & (\R.curInst\(20)))))) # (\R.curInst\(22) & ((((\Mux109~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (((\RegFile[2][13]~q\)))) 
-- # (\R.curInst\(20) & (\RegFile[3][13]~q\)))) # (\R.curInst\(22) & ((((\Mux109~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001010000010100010001001010101010111110101111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[3][13]~q\,
	datac => \ALT_INV_RegFile[2][13]~q\,
	datad => \ALT_INV_R.curInst\(20),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux109~0_combout\,
	datag => \ALT_INV_RegFile[1][13]~q\,
	combout => \Mux109~26_combout\);

-- Location: FF_X72_Y1_N8
\RegFile[23][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(13),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][13]~q\);

-- Location: FF_X71_Y1_N28
\RegFile[22][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(13),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][13]~q\);

-- Location: FF_X71_Y2_N14
\RegFile[21][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(13),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][13]~q\);

-- Location: FF_X72_Y1_N2
\RegFile[17][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(13),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][13]~q\);

-- Location: LABCELL_X73_Y1_N24
\RegFile[18][13]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[18][13]~feeder_combout\ = ( \R.regWriteData\(13) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(13),
	combout => \RegFile[18][13]~feeder_combout\);

-- Location: FF_X73_Y1_N25
\RegFile[18][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][13]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][13]~q\);

-- Location: FF_X72_Y1_N26
\RegFile[19][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(13),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][13]~q\);

-- Location: LABCELL_X77_Y2_N6
\RegFile[16][13]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[16][13]~feeder_combout\ = ( \R.regWriteData\(13) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(13),
	combout => \RegFile[16][13]~feeder_combout\);

-- Location: FF_X77_Y2_N7
\RegFile[16][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[16][13]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][13]~q\);

-- Location: MLABCELL_X72_Y1_N0
\Mux109~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux109~18_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[16][13]~q\))) # (\R.curInst\(20) & (\RegFile[17][13]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & (\RegFile[18][13]~q\)) # (\R.curInst\(20) & ((\RegFile[19][13]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[17][13]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[18][13]~q\,
	datad => \ALT_INV_RegFile[19][13]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][13]~q\,
	combout => \Mux109~18_combout\);

-- Location: FF_X71_Y1_N58
\RegFile[20][13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(13),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][13]~q\);

-- Location: LABCELL_X71_Y2_N12
\Mux109~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux109~5_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux109~18_combout\))))) # (\R.curInst\(22) & (((!\Mux109~18_combout\ & (\RegFile[20][13]~q\)) # (\Mux109~18_combout\ & ((\RegFile[21][13]~q\)))))) ) ) # ( \R.curInst\(21) & ( 
-- (!\R.curInst\(22) & ((((\Mux109~18_combout\))))) # (\R.curInst\(22) & (((!\Mux109~18_combout\ & ((\RegFile[22][13]~q\))) # (\Mux109~18_combout\ & (\RegFile[23][13]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110101010111111111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[23][13]~q\,
	datac => \ALT_INV_RegFile[22][13]~q\,
	datad => \ALT_INV_RegFile[21][13]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux109~18_combout\,
	datag => \ALT_INV_RegFile[20][13]~q\,
	combout => \Mux109~5_combout\);

-- Location: LABCELL_X71_Y2_N30
\Mux109~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux109~13_combout\ = ( \Mux109~26_combout\ & ( \Mux109~5_combout\ & ( (!\R.curInst\(23)) # ((!\R.curInst\(24) & ((\Mux109~1_combout\))) # (\R.curInst\(24) & (\Mux109~9_combout\))) ) ) ) # ( !\Mux109~26_combout\ & ( \Mux109~5_combout\ & ( 
-- (!\R.curInst\(23) & (\R.curInst\(24))) # (\R.curInst\(23) & ((!\R.curInst\(24) & ((\Mux109~1_combout\))) # (\R.curInst\(24) & (\Mux109~9_combout\)))) ) ) ) # ( \Mux109~26_combout\ & ( !\Mux109~5_combout\ & ( (!\R.curInst\(23) & (!\R.curInst\(24))) # 
-- (\R.curInst\(23) & ((!\R.curInst\(24) & ((\Mux109~1_combout\))) # (\R.curInst\(24) & (\Mux109~9_combout\)))) ) ) ) # ( !\Mux109~26_combout\ & ( !\Mux109~5_combout\ & ( (\R.curInst\(23) & ((!\R.curInst\(24) & ((\Mux109~1_combout\))) # (\R.curInst\(24) & 
-- (\Mux109~9_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000101000101100010011100110100100011011001111010101111101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(23),
	datab => \ALT_INV_R.curInst\(24),
	datac => \ALT_INV_Mux109~9_combout\,
	datad => \ALT_INV_Mux109~1_combout\,
	datae => \ALT_INV_Mux109~26_combout\,
	dataf => \ALT_INV_Mux109~5_combout\,
	combout => \Mux109~13_combout\);

-- Location: LABCELL_X71_Y6_N39
\NxR.aluData2[13]~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[13]~10_combout\ = ( \Mux109~13_combout\ & ( (!\vAluSrc2~1_combout\) # ((\Equal4~1_combout\ & \Mux141~0_combout\)) ) ) # ( !\Mux109~13_combout\ & ( (\Equal4~1_combout\ & (\Mux141~0_combout\ & \vAluSrc2~1_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000011000000000000001111111111000000111111111100000011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Equal4~1_combout\,
	datac => \ALT_INV_Mux141~0_combout\,
	datad => \ALT_INV_vAluSrc2~1_combout\,
	dataf => \ALT_INV_Mux109~13_combout\,
	combout => \NxR.aluData2[13]~10_combout\);

-- Location: FF_X71_Y6_N16
\R.aluData2[13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \NxR.aluData2[13]~10_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData2\(13));

-- Location: LABCELL_X79_Y8_N18
\vAluRes~56\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~56_combout\ = ( !\R.aluCalc~q\ & ( (((\R.aluRes\(13)))) ) ) # ( \R.aluCalc~q\ & ( ((!\Add1~53_sumout\ & (\Add2~53_sumout\ & ((\R.aluOp.ALUOpSub~q\)))) # (\Add1~53_sumout\ & (((\Add2~53_sumout\ & \R.aluOp.ALUOpSub~q\)) # (\R.aluOp.ALUOpAdd~q\)))) 
-- # (\Selector19~3_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100001111000001010011011100001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add1~53_sumout\,
	datab => \ALT_INV_Add2~53_sumout\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datae => \ALT_INV_R.aluCalc~q\,
	dataf => \ALT_INV_Selector19~3_combout\,
	datag => \ALT_INV_R.aluRes\(13),
	combout => \vAluRes~56_combout\);

-- Location: MLABCELL_X78_Y7_N42
\Comb:vJumpAdr[13]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[13]~0_combout\ = ( \Add3~53_sumout\ & ( (!\Equal4~2_combout\) # (\vAluRes~56_combout\) ) ) # ( !\Add3~53_sumout\ & ( (\vAluRes~56_combout\ & \Equal4~2_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000110000001111110011111100111111001111110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_vAluRes~56_combout\,
	datac => \ALT_INV_Equal4~2_combout\,
	dataf => \ALT_INV_Add3~53_sumout\,
	combout => \Comb:vJumpAdr[13]~0_combout\);

-- Location: FF_X78_Y7_N43
\R.curPC[13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[13]~0_combout\,
	asdata => \Add0~45_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(13));

-- Location: LABCELL_X70_Y2_N18
\Mux77~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux77~14_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[8][13]~q\))) # (\R.curInst\(15) & (\RegFile[9][13]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[10][13]~q\))) # (\R.curInst\(15) & (\RegFile[11][13]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[11][13]~q\,
	datab => \ALT_INV_RegFile[9][13]~q\,
	datac => \ALT_INV_RegFile[10][13]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][13]~q\,
	combout => \Mux77~14_combout\);

-- Location: LABCELL_X70_Y2_N24
\Mux77~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux77~1_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux77~14_combout\)))) # (\R.curInst\(17) & ((!\Mux77~14_combout\ & ((\RegFile[12][13]~q\))) # (\Mux77~14_combout\ & (\RegFile[13][13]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux77~14_combout\)))) # (\R.curInst\(17) & ((!\Mux77~14_combout\ & ((\RegFile[14][13]~q\))) # (\Mux77~14_combout\ & (\RegFile[15][13]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][13]~q\,
	datab => \ALT_INV_RegFile[15][13]~q\,
	datac => \ALT_INV_RegFile[14][13]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux77~14_combout\,
	datag => \ALT_INV_RegFile[12][13]~q\,
	combout => \Mux77~1_combout\);

-- Location: MLABCELL_X72_Y1_N24
\Mux77~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux77~18_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[16][13]~q\))) # (\R.curInst\(15) & (\RegFile[17][13]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & (\RegFile[18][13]~q\)) # (\R.curInst\(15) & ((\RegFile[19][13]~q\))))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[17][13]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[18][13]~q\,
	datad => \ALT_INV_RegFile[19][13]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][13]~q\,
	combout => \Mux77~18_combout\);

-- Location: MLABCELL_X72_Y1_N6
\Mux77~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux77~5_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux77~18_combout\))))) # (\R.curInst\(17) & (((!\Mux77~18_combout\ & (\RegFile[20][13]~q\)) # (\Mux77~18_combout\ & ((\RegFile[21][13]~q\)))))) ) ) # ( \R.curInst\(16) & ( 
-- (!\R.curInst\(17) & ((((\Mux77~18_combout\))))) # (\R.curInst\(17) & (((!\Mux77~18_combout\ & ((\RegFile[22][13]~q\))) # (\Mux77~18_combout\ & (\RegFile[23][13]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110101010111111111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[23][13]~q\,
	datac => \ALT_INV_RegFile[22][13]~q\,
	datad => \ALT_INV_RegFile[21][13]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux77~18_combout\,
	datag => \ALT_INV_RegFile[20][13]~q\,
	combout => \Mux77~5_combout\);

-- Location: LABCELL_X67_Y2_N18
\Mux77~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux77~22_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[24][13]~q\))) # (\R.curInst\(15) & (\RegFile[25][13]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[26][13]~q\))) # (\R.curInst\(15) & (\RegFile[27][13]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[27][13]~q\,
	datab => \ALT_INV_RegFile[25][13]~q\,
	datac => \ALT_INV_RegFile[26][13]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][13]~q\,
	combout => \Mux77~22_combout\);

-- Location: LABCELL_X73_Y2_N36
\Mux77~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux77~9_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux77~22_combout\)))) # (\R.curInst\(17) & ((!\Mux77~22_combout\ & ((\RegFile[28][13]~q\))) # (\Mux77~22_combout\ & (\RegFile[29][13]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux77~22_combout\)))) # (\R.curInst\(17) & ((!\Mux77~22_combout\ & ((\RegFile[30][13]~q\))) # (\Mux77~22_combout\ & (\RegFile[31][13]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][13]~q\,
	datab => \ALT_INV_RegFile[29][13]~q\,
	datac => \ALT_INV_RegFile[30][13]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux77~22_combout\,
	datag => \ALT_INV_RegFile[28][13]~q\,
	combout => \Mux77~9_combout\);

-- Location: LABCELL_X73_Y3_N42
\Mux77~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux77~0_combout\ = ( \RegFile[7][13]~q\ & ( \R.curInst\(15) & ( (\R.curInst\(16)) # (\RegFile[5][13]~q\) ) ) ) # ( !\RegFile[7][13]~q\ & ( \R.curInst\(15) & ( (\RegFile[5][13]~q\ & !\R.curInst\(16)) ) ) ) # ( \RegFile[7][13]~q\ & ( !\R.curInst\(15) & ( 
-- (!\R.curInst\(16) & (\RegFile[4][13]~q\)) # (\R.curInst\(16) & ((\RegFile[6][13]~q\))) ) ) ) # ( !\RegFile[7][13]~q\ & ( !\R.curInst\(15) & ( (!\R.curInst\(16) & (\RegFile[4][13]~q\)) # (\R.curInst\(16) & ((\RegFile[6][13]~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010100001111010101010000111100110011000000000011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[4][13]~q\,
	datab => \ALT_INV_RegFile[5][13]~q\,
	datac => \ALT_INV_RegFile[6][13]~q\,
	datad => \ALT_INV_R.curInst\(16),
	datae => \ALT_INV_RegFile[7][13]~q\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux77~0_combout\);

-- Location: LABCELL_X73_Y3_N6
\Mux77~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux77~26_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((\RegFile[1][13]~q\ & ((\R.curInst\(15))))))) # (\R.curInst\(17) & ((((\Mux77~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[2][13]~q\))) # 
-- (\R.curInst\(15) & (\RegFile[3][13]~q\))))) # (\R.curInst\(17) & ((((\Mux77~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000001010101000010100101111100001010010111110010001001110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[3][13]~q\,
	datac => \ALT_INV_RegFile[2][13]~q\,
	datad => \ALT_INV_Mux77~0_combout\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[1][13]~q\,
	combout => \Mux77~26_combout\);

-- Location: LABCELL_X73_Y2_N9
\Mux77~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux77~13_combout\ = ( \Mux77~9_combout\ & ( \Mux77~26_combout\ & ( (!\R.curInst\(18) & ((!\R.curInst\(19)) # ((\Mux77~5_combout\)))) # (\R.curInst\(18) & (((\Mux77~1_combout\)) # (\R.curInst\(19)))) ) ) ) # ( !\Mux77~9_combout\ & ( \Mux77~26_combout\ & ( 
-- (!\R.curInst\(18) & ((!\R.curInst\(19)) # ((\Mux77~5_combout\)))) # (\R.curInst\(18) & (!\R.curInst\(19) & (\Mux77~1_combout\))) ) ) ) # ( \Mux77~9_combout\ & ( !\Mux77~26_combout\ & ( (!\R.curInst\(18) & (\R.curInst\(19) & ((\Mux77~5_combout\)))) # 
-- (\R.curInst\(18) & (((\Mux77~1_combout\)) # (\R.curInst\(19)))) ) ) ) # ( !\Mux77~9_combout\ & ( !\Mux77~26_combout\ & ( (!\R.curInst\(18) & (\R.curInst\(19) & ((\Mux77~5_combout\)))) # (\R.curInst\(18) & (!\R.curInst\(19) & (\Mux77~1_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010000100110000101010011011110001100101011101001110110111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(18),
	datab => \ALT_INV_R.curInst\(19),
	datac => \ALT_INV_Mux77~1_combout\,
	datad => \ALT_INV_Mux77~5_combout\,
	datae => \ALT_INV_Mux77~9_combout\,
	dataf => \ALT_INV_Mux77~26_combout\,
	combout => \Mux77~13_combout\);

-- Location: LABCELL_X74_Y6_N12
\Mux241~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux241~0_combout\ = ( \Mux77~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC\(13)))) ) ) # ( !\Mux77~13_combout\ & ( (!\vAluSrc1~1_combout\ & (\vAluSrc1~2_combout\ & \R.curPC\(13))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001000000010000000100000001010001010100010101000101010001010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluSrc1~1_combout\,
	datab => \ALT_INV_vAluSrc1~2_combout\,
	datac => \ALT_INV_R.curPC\(13),
	dataf => \ALT_INV_Mux77~13_combout\,
	combout => \Mux241~0_combout\);

-- Location: LABCELL_X74_Y6_N30
\ShiftRight1~36\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~36_combout\ = ( \Mux242~0_combout\ & ( \Mux243~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\) # ((!\NxR.aluData2[0]~16_combout\ & ((\Mux241~0_combout\))) # (\NxR.aluData2[0]~16_combout\ & (\Mux240~0_combout\))) ) ) ) # ( !\Mux242~0_combout\ & 
-- ( \Mux243~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (((!\NxR.aluData2[1]~17_combout\) # (\Mux241~0_combout\)))) # (\NxR.aluData2[0]~16_combout\ & (\Mux240~0_combout\ & ((\NxR.aluData2[1]~17_combout\)))) ) ) ) # ( \Mux242~0_combout\ & ( 
-- !\Mux243~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (((\Mux241~0_combout\ & \NxR.aluData2[1]~17_combout\)))) # (\NxR.aluData2[0]~16_combout\ & (((!\NxR.aluData2[1]~17_combout\)) # (\Mux240~0_combout\))) ) ) ) # ( !\Mux242~0_combout\ & ( 
-- !\Mux243~0_combout\ & ( (\NxR.aluData2[1]~17_combout\ & ((!\NxR.aluData2[0]~16_combout\ & ((\Mux241~0_combout\))) # (\NxR.aluData2[0]~16_combout\ & (\Mux240~0_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110101000011110011010111110000001101011111111100110101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux240~0_combout\,
	datab => \ALT_INV_Mux241~0_combout\,
	datac => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datad => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datae => \ALT_INV_Mux242~0_combout\,
	dataf => \ALT_INV_Mux243~0_combout\,
	combout => \ShiftRight1~36_combout\);

-- Location: FF_X74_Y6_N31
\ShiftRight1~36_NEW_REG280\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~36_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~36_OTERM281\);

-- Location: LABCELL_X73_Y7_N6
\ShiftRight1~34\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~34_combout\ = ( \NxR.aluData2[0]~16_combout\ & ( \Mux250~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\) # (\Mux248~0_combout\) ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( \Mux250~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & 
-- ((\Mux251~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux249~0_combout\)) ) ) ) # ( \NxR.aluData2[0]~16_combout\ & ( !\Mux250~0_combout\ & ( (\Mux248~0_combout\ & \NxR.aluData2[1]~17_combout\) ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( 
-- !\Mux250~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((\Mux251~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux249~0_combout\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100110011000000000101010100001111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux248~0_combout\,
	datab => \ALT_INV_Mux249~0_combout\,
	datac => \ALT_INV_Mux251~0_combout\,
	datad => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datae => \ALT_INV_NxR.aluData2[0]~16_combout\,
	dataf => \ALT_INV_Mux250~0_combout\,
	combout => \ShiftRight1~34_combout\);

-- Location: FF_X73_Y7_N7
\ShiftRight1~38_OTERM439_NEW_REG744\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~34_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~38_OTERM439_OTERM745\);

-- Location: LABCELL_X77_Y7_N54
\ShiftRight1~38\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~38_combout\ = ( \ShiftRight1~38_OTERM439_OTERM745\ & ( \R.aluData2\(3) & ( (!\R.aluData2\(2) & (\ShiftRight1~36_OTERM281\)) # (\R.aluData2\(2) & ((\ShiftRight1~37_OTERM283\))) ) ) ) # ( !\ShiftRight1~38_OTERM439_OTERM745\ & ( \R.aluData2\(3) 
-- & ( (!\R.aluData2\(2) & (\ShiftRight1~36_OTERM281\)) # (\R.aluData2\(2) & ((\ShiftRight1~37_OTERM283\))) ) ) ) # ( \ShiftRight1~38_OTERM439_OTERM745\ & ( !\R.aluData2\(3) & ( (!\R.aluData2\(2)) # (\ShiftRight1~35_OTERM279\) ) ) ) # ( 
-- !\ShiftRight1~38_OTERM439_OTERM745\ & ( !\R.aluData2\(3) & ( (\ShiftRight1~35_OTERM279\ & \R.aluData2\(2)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110011111111110011001101010101000011110101010100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~36_OTERM281\,
	datab => \ALT_INV_ShiftRight1~35_OTERM279\,
	datac => \ALT_INV_ShiftRight1~37_OTERM283\,
	datad => \ALT_INV_R.aluData2\(2),
	datae => \ALT_INV_ShiftRight1~38_OTERM439_OTERM745\,
	dataf => \ALT_INV_R.aluData2\(3),
	combout => \ShiftRight1~38_combout\);

-- Location: MLABCELL_X82_Y7_N21
\Selector29~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector29~2_combout\ = ( \ShiftRight1~33_combout\ & ( (!\Selector31~6_OTERM381\ & (\Selector29~1_combout\ & ((!\Selector31~5_OTERM599\) # (!\ShiftRight1~38_combout\)))) ) ) # ( !\ShiftRight1~33_combout\ & ( (\Selector29~1_combout\ & 
-- ((!\Selector31~5_OTERM599\) # (!\ShiftRight1~38_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110000001100110011000000100010001000000010001000100000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector31~6_OTERM381\,
	datab => \ALT_INV_Selector29~1_combout\,
	datac => \ALT_INV_Selector31~5_OTERM599\,
	datad => \ALT_INV_ShiftRight1~38_combout\,
	dataf => \ALT_INV_ShiftRight1~33_combout\,
	combout => \Selector29~2_combout\);

-- Location: LABCELL_X83_Y6_N54
\Selector29~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector29~3_combout\ = ( \Add1~13_sumout\ & ( ((\R.aluOp.ALUOpSub~q\ & \Add2~13_sumout\)) # (\R.aluOp.ALUOpAdd~q\) ) ) # ( !\Add1~13_sumout\ & ( (\R.aluOp.ALUOpSub~q\ & \Add2~13_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110011000000000011001100001111001111110000111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_Add2~13_sumout\,
	dataf => \ALT_INV_Add1~13_sumout\,
	combout => \Selector29~3_combout\);

-- Location: LABCELL_X83_Y5_N0
\Selector29~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector29~4_combout\ = ( \Selector29~2_combout\ & ( ((\ShiftRight0~5_combout\ & \Selector31~7_OTERM383\)) # (\Selector29~3_combout\) ) ) # ( !\Selector29~2_combout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111111111111111111100001111001111110000111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_ShiftRight0~5_combout\,
	datac => \ALT_INV_Selector29~3_combout\,
	datad => \ALT_INV_Selector31~7_OTERM383\,
	dataf => \ALT_INV_Selector29~2_combout\,
	combout => \Selector29~4_combout\);

-- Location: FF_X83_Y5_N2
\R.aluRes[3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector29~4_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(3));

-- Location: MLABCELL_X82_Y7_N9
\vAluRes~3_RESYN1066\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~3_RESYN1066_BDD1067\ = (!\R.aluOp.ALUOpSub~q\ & (\ShiftRight0~5_combout\ & ((\Selector31~7_OTERM383\)))) # (\R.aluOp.ALUOpSub~q\ & (((\ShiftRight0~5_combout\ & \Selector31~7_OTERM383\)) # (\Add2~13_sumout\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100110111000001010011011100000101001101110000010100110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datab => \ALT_INV_ShiftRight0~5_combout\,
	datac => \ALT_INV_Add2~13_sumout\,
	datad => \ALT_INV_Selector31~7_OTERM383\,
	combout => \vAluRes~3_RESYN1066_BDD1067\);

-- Location: MLABCELL_X82_Y7_N0
\vAluRes~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~3_combout\ = ( \Add1~13_sumout\ & ( \R.aluOp.ALUOpAdd~q\ & ( (\R.aluRes\(3)) # (\R.aluCalc~q\) ) ) ) # ( !\Add1~13_sumout\ & ( \R.aluOp.ALUOpAdd~q\ & ( (!\R.aluCalc~q\ & (((\R.aluRes\(3))))) # (\R.aluCalc~q\ & ((!\Selector29~2_combout\) # 
-- ((\vAluRes~3_RESYN1066_BDD1067\)))) ) ) ) # ( \Add1~13_sumout\ & ( !\R.aluOp.ALUOpAdd~q\ & ( (!\R.aluCalc~q\ & (((\R.aluRes\(3))))) # (\R.aluCalc~q\ & ((!\Selector29~2_combout\) # ((\vAluRes~3_RESYN1066_BDD1067\)))) ) ) ) # ( !\Add1~13_sumout\ & ( 
-- !\R.aluOp.ALUOpAdd~q\ & ( (!\R.aluCalc~q\ & (((\R.aluRes\(3))))) # (\R.aluCalc~q\ & ((!\Selector29~2_combout\) # ((\vAluRes~3_RESYN1066_BDD1067\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010111000111111001011100011111100101110001111110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector29~2_combout\,
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_R.aluRes\(3),
	datad => \ALT_INV_vAluRes~3_RESYN1066_BDD1067\,
	datae => \ALT_INV_Add1~13_sumout\,
	dataf => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	combout => \vAluRes~3_combout\);

-- Location: MLABCELL_X82_Y4_N48
\Comb:vJumpAdr[3]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[3]~0_combout\ = ( \Equal4~2_combout\ & ( \Add3~13_sumout\ & ( \vAluRes~3_combout\ ) ) ) # ( !\Equal4~2_combout\ & ( \Add3~13_sumout\ ) ) # ( \Equal4~2_combout\ & ( !\Add3~13_sumout\ & ( \vAluRes~3_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000001100110011001111111111111111110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_vAluRes~3_combout\,
	datae => \ALT_INV_Equal4~2_combout\,
	dataf => \ALT_INV_Add3~13_sumout\,
	combout => \Comb:vJumpAdr[3]~0_combout\);

-- Location: FF_X82_Y4_N49
\R.curPC[3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[3]~0_combout\,
	asdata => \Add0~5_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(3));

-- Location: LABCELL_X83_Y6_N57
\R.regWriteData[3]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.regWriteData[3]~feeder_combout\ = \Add0~5_sumout\

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101010101010101010101010101010101010101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add0~5_sumout\,
	combout => \R.regWriteData[3]~feeder_combout\);

-- Location: IOIBUF_X89_Y20_N44
\avm_d_readdata[27]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(27),
	o => \avm_d_readdata[27]~input_o\);

-- Location: LABCELL_X83_Y5_N48
\Comb:vRegWriteData[3]~0_RESYN1084\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[3]~0_RESYN1084_BDD1085\ = ( \Mux222~0_combout\ & ( \R.memToReg~q\ ) ) # ( \Mux222~0_combout\ & ( !\R.memToReg~q\ & ( (!\R.aluCalc~q\ & (\R.aluRes\(3))) # (\R.aluCalc~q\ & (((\Selector31~7_OTERM383\ & \ShiftRight0~5_combout\)))) ) ) ) # 
-- ( !\Mux222~0_combout\ & ( !\R.memToReg~q\ & ( (!\R.aluCalc~q\ & (\R.aluRes\(3))) # (\R.aluCalc~q\ & (((\Selector31~7_OTERM383\ & \ShiftRight0~5_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101000001010011010100000101001100000000000000001111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluRes\(3),
	datab => \ALT_INV_Selector31~7_OTERM383\,
	datac => \ALT_INV_R.aluCalc~q\,
	datad => \ALT_INV_ShiftRight0~5_combout\,
	datae => \ALT_INV_Mux222~0_combout\,
	dataf => \ALT_INV_R.memToReg~q\,
	combout => \Comb:vRegWriteData[3]~0_RESYN1084_BDD1085\);

-- Location: LABCELL_X83_Y6_N36
\Comb:vRegWriteData[3]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[3]~0_combout\ = ( \Selector29~3_combout\ & ( \Comb:vRegWriteData[3]~0_RESYN1084_BDD1085\ & ( (!\R.memToReg~q\) # (\avm_d_readdata[27]~input_o\) ) ) ) # ( !\Selector29~3_combout\ & ( \Comb:vRegWriteData[3]~0_RESYN1084_BDD1085\ & ( 
-- (!\R.memToReg~q\) # (\avm_d_readdata[27]~input_o\) ) ) ) # ( \Selector29~3_combout\ & ( !\Comb:vRegWriteData[3]~0_RESYN1084_BDD1085\ & ( (\R.aluCalc~q\ & !\R.memToReg~q\) ) ) ) # ( !\Selector29~3_combout\ & ( !\Comb:vRegWriteData[3]~0_RESYN1084_BDD1085\ & 
-- ( (!\Selector29~2_combout\ & (\R.aluCalc~q\ & !\R.memToReg~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010000000100000001100000011000011110000111111111111000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector29~2_combout\,
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_R.memToReg~q\,
	datad => \ALT_INV_avm_d_readdata[27]~input_o\,
	datae => \ALT_INV_Selector29~3_combout\,
	dataf => \ALT_INV_Comb:vRegWriteData[3]~0_RESYN1084_BDD1085\,
	combout => \Comb:vRegWriteData[3]~0_combout\);

-- Location: FF_X83_Y6_N59
\R.regWriteData[3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \R.regWriteData[3]~feeder_combout\,
	asdata => \Comb:vRegWriteData[3]~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(3));

-- Location: FF_X65_Y1_N32
\RegFile[13][3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(3),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][3]~q\);

-- Location: LABCELL_X66_Y1_N24
\Mux119~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux119~14_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[8][3]~q\))) # (\R.curInst\(20) & (\RegFile[9][3]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[10][3]~q\))) # (\R.curInst\(20) & (\RegFile[11][3]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][3]~q\,
	datab => \ALT_INV_RegFile[11][3]~q\,
	datac => \ALT_INV_RegFile[10][3]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][3]~q\,
	combout => \Mux119~14_combout\);

-- Location: LABCELL_X66_Y1_N39
\Mux119~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux119~1_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux119~14_combout\)))) # (\R.curInst\(22) & ((!\Mux119~14_combout\ & ((\RegFile[12][3]~q\))) # (\Mux119~14_combout\ & (\RegFile[13][3]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux119~14_combout\)))) # (\R.curInst\(22) & ((!\Mux119~14_combout\ & ((\RegFile[14][3]~q\))) # (\Mux119~14_combout\ & (\RegFile[15][3]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][3]~q\,
	datab => \ALT_INV_RegFile[15][3]~q\,
	datac => \ALT_INV_RegFile[14][3]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux119~14_combout\,
	datag => \ALT_INV_RegFile[12][3]~q\,
	combout => \Mux119~1_combout\);

-- Location: MLABCELL_X65_Y4_N42
\Mux119~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux119~22_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & (\RegFile[24][3]~q\)) # (\R.curInst\(20) & ((\RegFile[25][3]~q\)))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & ((\RegFile[26][3]~q\))) # (\R.curInst\(20) & (\RegFile[27][3]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001010101111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[27][3]~q\,
	datac => \ALT_INV_RegFile[26][3]~q\,
	datad => \ALT_INV_RegFile[25][3]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][3]~q\,
	combout => \Mux119~22_combout\);

-- Location: LABCELL_X68_Y6_N12
\Mux119~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux119~9_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux119~22_combout\)))) # (\R.curInst\(22) & ((!\Mux119~22_combout\ & ((\RegFile[28][3]~q\))) # (\Mux119~22_combout\ & (\RegFile[29][3]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux119~22_combout\)))) # (\R.curInst\(22) & ((!\Mux119~22_combout\ & ((\RegFile[30][3]~q\))) # (\Mux119~22_combout\ & (\RegFile[31][3]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[29][3]~q\,
	datab => \ALT_INV_RegFile[31][3]~q\,
	datac => \ALT_INV_RegFile[30][3]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux119~22_combout\,
	datag => \ALT_INV_RegFile[28][3]~q\,
	combout => \Mux119~9_combout\);

-- Location: LABCELL_X70_Y7_N42
\Mux119~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux119~18_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[16][3]~q\))) # (\R.curInst\(20) & (\RegFile[17][3]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & (\RegFile[18][3]~q\)) # (\R.curInst\(20) & ((\RegFile[19][3]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[17][3]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[18][3]~q\,
	datad => \ALT_INV_RegFile[19][3]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][3]~q\,
	combout => \Mux119~18_combout\);

-- Location: LABCELL_X70_Y7_N39
\Mux119~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux119~5_combout\ = ( !\R.curInst\(21) & ( ((!\Mux119~18_combout\ & (\RegFile[20][3]~q\ & (\R.curInst\(22)))) # (\Mux119~18_combout\ & (((!\R.curInst\(22)) # (\RegFile[21][3]~q\))))) ) ) # ( \R.curInst\(21) & ( (!\Mux119~18_combout\ & 
-- (((\RegFile[22][3]~q\ & (\R.curInst\(22)))))) # (\Mux119~18_combout\ & ((((!\R.curInst\(22)))) # (\RegFile[23][3]~q\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0011001100001100001100110001110100110011001111110011001100011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[23][3]~q\,
	datab => \ALT_INV_Mux119~18_combout\,
	datac => \ALT_INV_RegFile[22][3]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_RegFile[21][3]~q\,
	datag => \ALT_INV_RegFile[20][3]~q\,
	combout => \Mux119~5_combout\);

-- Location: LABCELL_X68_Y4_N42
\Mux119~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux119~0_combout\ = ( \RegFile[6][3]~q\ & ( \R.curInst\(21) & ( (!\R.curInst\(20)) # (\RegFile[7][3]~q\) ) ) ) # ( !\RegFile[6][3]~q\ & ( \R.curInst\(21) & ( (\RegFile[7][3]~q\ & \R.curInst\(20)) ) ) ) # ( \RegFile[6][3]~q\ & ( !\R.curInst\(21) & ( 
-- (!\R.curInst\(20) & ((\RegFile[4][3]~q\))) # (\R.curInst\(20) & (\RegFile[5][3]~q\)) ) ) ) # ( !\RegFile[6][3]~q\ & ( !\R.curInst\(21) & ( (!\R.curInst\(20) & ((\RegFile[4][3]~q\))) # (\R.curInst\(20) & (\RegFile[5][3]~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001101010101001100110101010100000000000011111111111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[5][3]~q\,
	datab => \ALT_INV_RegFile[4][3]~q\,
	datac => \ALT_INV_RegFile[7][3]~q\,
	datad => \ALT_INV_R.curInst\(20),
	datae => \ALT_INV_RegFile[6][3]~q\,
	dataf => \ALT_INV_R.curInst\(21),
	combout => \Mux119~0_combout\);

-- Location: LABCELL_X70_Y7_N24
\Mux119~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux119~26_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (\R.curInst\(20) & (((\RegFile[1][3]~q\))))) # (\R.curInst\(22) & (((\Mux119~0_combout\)))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (((\RegFile[2][3]~q\)))) # 
-- (\R.curInst\(20) & (((\RegFile[3][3]~q\)))))) # (\R.curInst\(22) & (((\Mux119~0_combout\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100110011000010100011001100000101001100110101111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(20),
	datab => \ALT_INV_Mux119~0_combout\,
	datac => \ALT_INV_RegFile[2][3]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_RegFile[3][3]~q\,
	datag => \ALT_INV_RegFile[1][3]~q\,
	combout => \Mux119~26_combout\);

-- Location: LABCELL_X70_Y7_N18
\Mux119~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux119~13_combout\ = ( \Mux119~5_combout\ & ( \Mux119~26_combout\ & ( (!\R.curInst\(23)) # ((!\R.curInst\(24) & (\Mux119~1_combout\)) # (\R.curInst\(24) & ((\Mux119~9_combout\)))) ) ) ) # ( !\Mux119~5_combout\ & ( \Mux119~26_combout\ & ( 
-- (!\R.curInst\(23) & (((!\R.curInst\(24))))) # (\R.curInst\(23) & ((!\R.curInst\(24) & (\Mux119~1_combout\)) # (\R.curInst\(24) & ((\Mux119~9_combout\))))) ) ) ) # ( \Mux119~5_combout\ & ( !\Mux119~26_combout\ & ( (!\R.curInst\(23) & (((\R.curInst\(24))))) 
-- # (\R.curInst\(23) & ((!\R.curInst\(24) & (\Mux119~1_combout\)) # (\R.curInst\(24) & ((\Mux119~9_combout\))))) ) ) ) # ( !\Mux119~5_combout\ & ( !\Mux119~26_combout\ & ( (\R.curInst\(23) & ((!\R.curInst\(24) & (\Mux119~1_combout\)) # (\R.curInst\(24) & 
-- ((\Mux119~9_combout\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100000101000100011010111110111011000001011011101110101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(23),
	datab => \ALT_INV_Mux119~1_combout\,
	datac => \ALT_INV_Mux119~9_combout\,
	datad => \ALT_INV_R.curInst\(24),
	datae => \ALT_INV_Mux119~5_combout\,
	dataf => \ALT_INV_Mux119~26_combout\,
	combout => \Mux119~13_combout\);

-- Location: LABCELL_X71_Y7_N3
\NxR.aluData2[3]~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[3]~18_combout\ = ( \Mux119~13_combout\ & ( (!\vAluSrc2~1_combout\) # ((\Equal4~1_combout\ & \Mux151~0_combout\)) ) ) # ( !\Mux119~13_combout\ & ( (\Equal4~1_combout\ & (\vAluSrc2~1_combout\ & \Mux151~0_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000101000000000000010111110000111101011111000011110101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Equal4~1_combout\,
	datac => \ALT_INV_vAluSrc2~1_combout\,
	datad => \ALT_INV_Mux151~0_combout\,
	dataf => \ALT_INV_Mux119~13_combout\,
	combout => \NxR.aluData2[3]~18_combout\);

-- Location: FF_X71_Y7_N16
\R.aluData2[3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \NxR.aluData2[3]~18_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData2\(3));

-- Location: LABCELL_X75_Y5_N24
\Selector7~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector7~2_combout\ = ( \R.aluData1\(25) & ( \R.aluData2[25]~DUPLICATE_q\ & ( ((\Selector17~0_OTERM391\) # (\R.aluOp.ALUOpOr~q\)) # (\R.aluOp.ALUOpAnd~DUPLICATE_q\) ) ) ) # ( !\R.aluData1\(25) & ( \R.aluData2[25]~DUPLICATE_q\ & ( 
-- ((\Selector17~0_OTERM391\) # (\R.aluOp.ALUOpOr~q\)) # (\R.aluOp.ALUOpXor~DUPLICATE_q\) ) ) ) # ( \R.aluData1\(25) & ( !\R.aluData2[25]~DUPLICATE_q\ & ( ((\Selector17~0_OTERM391\) # (\R.aluOp.ALUOpOr~q\)) # (\R.aluOp.ALUOpXor~DUPLICATE_q\) ) ) ) # ( 
-- !\R.aluData1\(25) & ( !\R.aluData2[25]~DUPLICATE_q\ & ( \Selector17~0_OTERM391\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111001111111111111100111111111111110101111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpAnd~DUPLICATE_q\,
	datab => \ALT_INV_R.aluOp.ALUOpXor~DUPLICATE_q\,
	datac => \ALT_INV_R.aluOp.ALUOpOr~q\,
	datad => \ALT_INV_Selector17~0_OTERM391\,
	datae => \ALT_INV_R.aluData1\(25),
	dataf => \ALT_INV_R.aluData2[25]~DUPLICATE_q\,
	combout => \Selector7~2_combout\);

-- Location: LABCELL_X75_Y5_N48
\Selector7~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector7~5_combout\ = ( !\R.aluData2\(2) & ( ((\Selector12~2_OTERM395\ & ((!\R.aluData2\(3) & ((\ShiftLeft0~12_OTERM791\))) # (\R.aluData2\(3) & (\ShiftLeft0~1_OTERM255\))))) # (\Selector7~2_combout\) ) ) # ( \R.aluData2\(2) & ( (((!\R.aluData2\(3) & 
-- (\Selector12~2_OTERM395\ & \ShiftLeft0~7_OTERM205\))) # (\Selector7~2_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000100100011000000100000001011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(3),
	datab => \ALT_INV_Selector12~2_OTERM395\,
	datac => \ALT_INV_ShiftLeft0~7_OTERM205\,
	datad => \ALT_INV_ShiftLeft0~12_OTERM791\,
	datae => \ALT_INV_R.aluData2\(2),
	dataf => \ALT_INV_Selector7~2_combout\,
	datag => \ALT_INV_ShiftLeft0~1_OTERM255\,
	combout => \Selector7~5_combout\);

-- Location: MLABCELL_X82_Y5_N39
\Selector7~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector7~4_combout\ = (!\Selector7~5_combout\ & !\Selector7~1_combout\)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111000000000000111100000000000011110000000000001111000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Selector7~5_combout\,
	datad => \ALT_INV_Selector7~1_combout\,
	combout => \Selector7~4_combout\);

-- Location: LABCELL_X79_Y5_N51
\vAluRes~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~25_combout\ = ( \Add1~101_sumout\ & ( \Add2~101_sumout\ & ( (\R.aluCalc~q\ & (((!\Selector7~4_combout\) # (\R.aluOp.ALUOpAdd~q\)) # (\R.aluOp.ALUOpSub~q\))) ) ) ) # ( !\Add1~101_sumout\ & ( \Add2~101_sumout\ & ( (\R.aluCalc~q\ & 
-- ((!\Selector7~4_combout\) # (\R.aluOp.ALUOpSub~q\))) ) ) ) # ( \Add1~101_sumout\ & ( !\Add2~101_sumout\ & ( (\R.aluCalc~q\ & ((!\Selector7~4_combout\) # (\R.aluOp.ALUOpAdd~q\))) ) ) ) # ( !\Add1~101_sumout\ & ( !\Add2~101_sumout\ & ( 
-- (!\Selector7~4_combout\ & \R.aluCalc~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011001100000000001100111100000000110111010000000011011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datab => \ALT_INV_Selector7~4_combout\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_R.aluCalc~q\,
	datae => \ALT_INV_Add1~101_sumout\,
	dataf => \ALT_INV_Add2~101_sumout\,
	combout => \vAluRes~25_combout\);

-- Location: MLABCELL_X78_Y4_N24
\Comb:vJumpAdr[25]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[25]~0_combout\ = ( \Add3~101_sumout\ & ( (!\Equal4~2_combout\) # ((\vAluRes~26_combout\) # (\vAluRes~25_combout\)) ) ) # ( !\Add3~101_sumout\ & ( (\Equal4~2_combout\ & ((\vAluRes~26_combout\) # (\vAluRes~25_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001010100010101000101010001010110111111101111111011111110111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Equal4~2_combout\,
	datab => \ALT_INV_vAluRes~25_combout\,
	datac => \ALT_INV_vAluRes~26_combout\,
	dataf => \ALT_INV_Add3~101_sumout\,
	combout => \Comb:vJumpAdr[25]~0_combout\);

-- Location: FF_X78_Y4_N25
\R.curPC[25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[25]~0_combout\,
	asdata => \Add0~93_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(25));

-- Location: LABCELL_X81_Y5_N42
\Add0~97\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~97_sumout\ = SUM(( \R.curPC\(26) ) + ( GND ) + ( \Add0~94\ ))
-- \Add0~98\ = CARRY(( \R.curPC\(26) ) + ( GND ) + ( \Add0~94\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.curPC\(26),
	cin => \Add0~94\,
	sumout => \Add0~97_sumout\,
	cout => \Add0~98\);

-- Location: IOIBUF_X36_Y81_N18
\avm_d_readdata[2]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(2),
	o => \avm_d_readdata[2]~input_o\);

-- Location: LABCELL_X79_Y2_N9
\Comb:vRegWriteData[26]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[26]~1_combout\ = ( \avm_d_readdata[23]~input_o\ & ( \avm_d_readdata[2]~input_o\ & ( (!\R.curInst\(14) & ((!\R.curInst\(12) & ((\R.curInst\(13)) # (\avm_d_readdata[31]~input_o\))) # (\R.curInst\(12) & ((!\R.curInst\(13)))))) ) ) ) # ( 
-- !\avm_d_readdata[23]~input_o\ & ( \avm_d_readdata[2]~input_o\ & ( (!\R.curInst\(12) & (!\R.curInst\(14) & ((\R.curInst\(13)) # (\avm_d_readdata[31]~input_o\)))) ) ) ) # ( \avm_d_readdata[23]~input_o\ & ( !\avm_d_readdata[2]~input_o\ & ( (!\R.curInst\(14) 
-- & (!\R.curInst\(13) & ((\avm_d_readdata[31]~input_o\) # (\R.curInst\(12))))) ) ) ) # ( !\avm_d_readdata[23]~input_o\ & ( !\avm_d_readdata[2]~input_o\ & ( (!\R.curInst\(12) & (\avm_d_readdata[31]~input_o\ & (!\R.curInst\(14) & !\R.curInst\(13)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010000000000000011100000000000000100000101000000111000010100000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(12),
	datab => \ALT_INV_avm_d_readdata[31]~input_o\,
	datac => \ALT_INV_R.curInst\(14),
	datad => \ALT_INV_R.curInst\(13),
	datae => \ALT_INV_avm_d_readdata[23]~input_o\,
	dataf => \ALT_INV_avm_d_readdata[2]~input_o\,
	combout => \Comb:vRegWriteData[26]~1_combout\);

-- Location: MLABCELL_X78_Y7_N12
\Comb:vRegWriteData[26]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[26]~2_combout\ = ( \Comb:vRegWriteData[26]~1_combout\ & ( (\Selector6~1_combout\ & (!\R.memToReg~q\ & ((!\Add1~105_sumout\) # (!\R.aluOp.ALUOpAdd~q\)))) ) ) # ( !\Comb:vRegWriteData[26]~1_combout\ & ( ((\Selector6~1_combout\ & 
-- ((!\Add1~105_sumout\) # (!\R.aluOp.ALUOpAdd~q\)))) # (\R.memToReg~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101111101001111010111110100111101010000010000000101000001000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector6~1_combout\,
	datab => \ALT_INV_Add1~105_sumout\,
	datac => \ALT_INV_R.memToReg~q\,
	datad => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	dataf => \ALT_INV_Comb:vRegWriteData[26]~1_combout\,
	combout => \Comb:vRegWriteData[26]~2_combout\);

-- Location: MLABCELL_X78_Y7_N18
\Comb:vRegWriteData[26]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[26]~0_combout\ = ( \Add2~105_sumout\ & ( \Comb:vRegWriteData[26]~2_combout\ & ( (!\R.memToReg~q\ & ((!\R.aluCalc~q\ & (\R.aluRes\(26))) # (\R.aluCalc~q\ & ((\R.aluOp.ALUOpSub~q\))))) ) ) ) # ( !\Add2~105_sumout\ & ( 
-- \Comb:vRegWriteData[26]~2_combout\ & ( (!\R.memToReg~q\ & (\R.aluRes\(26) & !\R.aluCalc~q\)) ) ) ) # ( \Add2~105_sumout\ & ( !\Comb:vRegWriteData[26]~2_combout\ & ( ((\R.aluCalc~q\) # (\R.aluRes\(26))) # (\R.memToReg~q\) ) ) ) # ( !\Add2~105_sumout\ & ( 
-- !\Comb:vRegWriteData[26]~2_combout\ & ( ((\R.aluCalc~q\) # (\R.aluRes\(26))) # (\R.memToReg~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0111011111111111011101111111111100100010000000000010001000001010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.memToReg~q\,
	datab => \ALT_INV_R.aluRes\(26),
	datac => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datad => \ALT_INV_R.aluCalc~q\,
	datae => \ALT_INV_Add2~105_sumout\,
	dataf => \ALT_INV_Comb:vRegWriteData[26]~2_combout\,
	combout => \Comb:vRegWriteData[26]~0_combout\);

-- Location: FF_X81_Y5_N44
\R.regWriteData[26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Add0~97_sumout\,
	asdata => \Comb:vRegWriteData[26]~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(26));

-- Location: FF_X70_Y6_N44
\RegFile[21][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(26),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][26]~q\);

-- Location: LABCELL_X70_Y4_N6
\Mux64~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux64~18_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & (\RegFile[16][26]~q\)) # (\R.curInst\(15) & ((\RegFile[17][26]~q\)))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & ((\RegFile[18][26]~q\))) # (\R.curInst\(15) & (\RegFile[19][26]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001010101111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[19][26]~q\,
	datac => \ALT_INV_RegFile[18][26]~q\,
	datad => \ALT_INV_RegFile[17][26]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][26]~q\,
	combout => \Mux64~18_combout\);

-- Location: LABCELL_X73_Y4_N24
\Mux64~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux64~5_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux64~18_combout\))))) # (\R.curInst\(17) & (((!\Mux64~18_combout\ & ((\RegFile[20][26]~q\))) # (\Mux64~18_combout\ & (\RegFile[21][26]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux64~18_combout\)))) # (\R.curInst\(17) & ((!\Mux64~18_combout\ & (\RegFile[22][26]~q\)) # (\Mux64~18_combout\ & ((\RegFile[23][26]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][26]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[22][26]~q\,
	datad => \ALT_INV_RegFile[23][26]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux64~18_combout\,
	datag => \ALT_INV_RegFile[20][26]~q\,
	combout => \Mux64~5_combout\);

-- Location: FF_X60_Y4_N40
\RegFile[2][26]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(26),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][26]~DUPLICATE_q\);

-- Location: FF_X61_Y4_N50
\RegFile[7][26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(26),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][26]~q\);

-- Location: LABCELL_X61_Y4_N12
\Mux64~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux64~0_combout\ = ( \R.curInst\(16) & ( \R.curInst\(15) & ( \RegFile[7][26]~q\ ) ) ) # ( !\R.curInst\(16) & ( \R.curInst\(15) & ( \RegFile[5][26]~q\ ) ) ) # ( \R.curInst\(16) & ( !\R.curInst\(15) & ( \RegFile[6][26]~q\ ) ) ) # ( !\R.curInst\(16) & ( 
-- !\R.curInst\(15) & ( \RegFile[4][26]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111001100110011001100000000111111110101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[7][26]~q\,
	datab => \ALT_INV_RegFile[6][26]~q\,
	datac => \ALT_INV_RegFile[4][26]~q\,
	datad => \ALT_INV_RegFile[5][26]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux64~0_combout\);

-- Location: LABCELL_X61_Y4_N24
\Mux64~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux64~26_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (\RegFile[1][26]~q\ & (\R.curInst\(15)))) # (\R.curInst\(17) & (((\Mux64~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & ((!\R.curInst\(15) & 
-- (((\RegFile[2][26]~DUPLICATE_q\)))) # (\R.curInst\(15) & (\RegFile[3][26]~q\)))) # (\R.curInst\(17) & ((((\Mux64~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001100000011000100010000110011001111110011111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][26]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[2][26]~DUPLICATE_q\,
	datad => \ALT_INV_R.curInst\(15),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux64~0_combout\,
	datag => \ALT_INV_RegFile[1][26]~q\,
	combout => \Mux64~26_combout\);

-- Location: LABCELL_X67_Y4_N42
\Mux64~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux64~22_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[24][26]~q\))) # (\R.curInst\(15) & (\RegFile[25][26]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & (\RegFile[26][26]~q\)) # (\R.curInst\(15) & ((\RegFile[27][26]~q\))))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[25][26]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[26][26]~q\,
	datad => \ALT_INV_RegFile[27][26]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][26]~q\,
	combout => \Mux64~22_combout\);

-- Location: LABCELL_X73_Y4_N54
\Mux64~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux64~9_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux64~22_combout\))))) # (\R.curInst\(17) & (((!\Mux64~22_combout\ & ((\RegFile[28][26]~q\))) # (\Mux64~22_combout\ & (\RegFile[29][26]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux64~22_combout\)))) # (\R.curInst\(17) & ((!\Mux64~22_combout\ & (\RegFile[30][26]~q\)) # (\Mux64~22_combout\ & ((\RegFile[31][26]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[29][26]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[30][26]~q\,
	datad => \ALT_INV_RegFile[31][26]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux64~22_combout\,
	datag => \ALT_INV_RegFile[28][26]~q\,
	combout => \Mux64~9_combout\);

-- Location: FF_X64_Y8_N32
\RegFile[10][26]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(26),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][26]~DUPLICATE_q\);

-- Location: LABCELL_X63_Y8_N6
\Mux64~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux64~14_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[8][26]~q\))) # (\R.curInst\(15) & (\RegFile[9][26]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & (\RegFile[10][26]~DUPLICATE_q\)) # (\R.curInst\(15) & ((\RegFile[11][26]~q\))))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][26]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[10][26]~DUPLICATE_q\,
	datad => \ALT_INV_RegFile[11][26]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][26]~q\,
	combout => \Mux64~14_combout\);

-- Location: LABCELL_X63_Y8_N18
\Mux64~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux64~1_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux64~14_combout\)))) # (\R.curInst\(17) & ((!\Mux64~14_combout\ & ((\RegFile[12][26]~q\))) # (\Mux64~14_combout\ & (\RegFile[13][26]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux64~14_combout\)))) # (\R.curInst\(17) & ((!\Mux64~14_combout\ & ((\RegFile[14][26]~q\))) # (\Mux64~14_combout\ & (\RegFile[15][26]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][26]~q\,
	datab => \ALT_INV_RegFile[13][26]~q\,
	datac => \ALT_INV_RegFile[14][26]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux64~14_combout\,
	datag => \ALT_INV_RegFile[12][26]~q\,
	combout => \Mux64~1_combout\);

-- Location: LABCELL_X73_Y4_N6
\Mux64~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux64~13_combout\ = ( \Mux64~9_combout\ & ( \Mux64~1_combout\ & ( ((!\R.curInst\(19) & ((\Mux64~26_combout\))) # (\R.curInst\(19) & (\Mux64~5_combout\))) # (\R.curInst\(18)) ) ) ) # ( !\Mux64~9_combout\ & ( \Mux64~1_combout\ & ( (!\R.curInst\(18) & 
-- ((!\R.curInst\(19) & ((\Mux64~26_combout\))) # (\R.curInst\(19) & (\Mux64~5_combout\)))) # (\R.curInst\(18) & (((!\R.curInst\(19))))) ) ) ) # ( \Mux64~9_combout\ & ( !\Mux64~1_combout\ & ( (!\R.curInst\(18) & ((!\R.curInst\(19) & ((\Mux64~26_combout\))) # 
-- (\R.curInst\(19) & (\Mux64~5_combout\)))) # (\R.curInst\(18) & (((\R.curInst\(19))))) ) ) ) # ( !\Mux64~9_combout\ & ( !\Mux64~1_combout\ & ( (!\R.curInst\(18) & ((!\R.curInst\(19) & ((\Mux64~26_combout\))) # (\R.curInst\(19) & (\Mux64~5_combout\)))) ) ) 
-- )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010011000100000001111100011100110100111101000011011111110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux64~5_combout\,
	datab => \ALT_INV_R.curInst\(18),
	datac => \ALT_INV_R.curInst\(19),
	datad => \ALT_INV_Mux64~26_combout\,
	datae => \ALT_INV_Mux64~9_combout\,
	dataf => \ALT_INV_Mux64~1_combout\,
	combout => \Mux64~13_combout\);

-- Location: LABCELL_X73_Y4_N42
\Mux228~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux228~0_combout\ = ( \Mux64~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC\(26)))) ) ) # ( !\Mux64~13_combout\ & ( (\vAluSrc1~2_combout\ & (!\vAluSrc1~1_combout\ & \R.curPC\(26))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010000000100000001000000010010001100100011001000110010001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluSrc1~2_combout\,
	datab => \ALT_INV_vAluSrc1~1_combout\,
	datac => \ALT_INV_R.curPC\(26),
	dataf => \ALT_INV_Mux64~13_combout\,
	combout => \Mux228~0_combout\);

-- Location: LABCELL_X73_Y4_N36
\ShiftRight1~12\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~12_combout\ = ( \Mux226~0_combout\ & ( \Mux227~0_combout\ & ( ((!\NxR.aluData2[0]~16_combout\ & ((\Mux229~0_combout\))) # (\NxR.aluData2[0]~16_combout\ & (\Mux228~0_combout\))) # (\NxR.aluData2[1]~17_combout\) ) ) ) # ( !\Mux226~0_combout\ & 
-- ( \Mux227~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (((\Mux229~0_combout\) # (\NxR.aluData2[1]~17_combout\)))) # (\NxR.aluData2[0]~16_combout\ & (\Mux228~0_combout\ & (!\NxR.aluData2[1]~17_combout\))) ) ) ) # ( \Mux226~0_combout\ & ( 
-- !\Mux227~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (((!\NxR.aluData2[1]~17_combout\ & \Mux229~0_combout\)))) # (\NxR.aluData2[0]~16_combout\ & (((\NxR.aluData2[1]~17_combout\)) # (\Mux228~0_combout\))) ) ) ) # ( !\Mux226~0_combout\ & ( 
-- !\Mux227~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((!\NxR.aluData2[0]~16_combout\ & ((\Mux229~0_combout\))) # (\NxR.aluData2[0]~16_combout\ & (\Mux228~0_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000010110000000101011011010100011010101110100001111110111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datab => \ALT_INV_Mux228~0_combout\,
	datac => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datad => \ALT_INV_Mux229~0_combout\,
	datae => \ALT_INV_Mux226~0_combout\,
	dataf => \ALT_INV_Mux227~0_combout\,
	combout => \ShiftRight1~12_combout\);

-- Location: FF_X73_Y4_N37
\ShiftRight1~12_NEW_REG56\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~12_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~12_OTERM57\);

-- Location: LABCELL_X77_Y9_N3
\ShiftRight0~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight0~1_combout\ = ( \R.aluData2\(3) & ( \ShiftRight0~0_OTERM17\ & ( (\R.aluData2\(2)) # (\ShiftRight1~12_OTERM57\) ) ) ) # ( !\R.aluData2\(3) & ( \ShiftRight0~0_OTERM17\ & ( (!\R.aluData2\(2) & ((\ShiftRight1~10_OTERM265\))) # (\R.aluData2\(2) & 
-- (\ShiftRight1~11_OTERM35\)) ) ) ) # ( \R.aluData2\(3) & ( !\ShiftRight0~0_OTERM17\ & ( (\ShiftRight1~12_OTERM57\ & !\R.aluData2\(2)) ) ) ) # ( !\R.aluData2\(3) & ( !\ShiftRight0~0_OTERM17\ & ( (!\R.aluData2\(2) & ((\ShiftRight1~10_OTERM265\))) # 
-- (\R.aluData2\(2) & (\ShiftRight1~11_OTERM35\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001111001111010001000100010000000011110011110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~12_OTERM57\,
	datab => \ALT_INV_R.aluData2\(2),
	datac => \ALT_INV_ShiftRight1~11_OTERM35\,
	datad => \ALT_INV_ShiftRight1~10_OTERM265\,
	datae => \ALT_INV_R.aluData2\(3),
	dataf => \ALT_INV_ShiftRight0~0_OTERM17\,
	combout => \ShiftRight0~1_combout\);

-- Location: MLABCELL_X72_Y7_N6
\ShiftRight1~15\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~15_combout\ = ( \NxR.aluData2[0]~16_combout\ & ( \Mux253~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((\Mux252~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & (\Mux250~0_combout\)) ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( 
-- \Mux253~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\) # (\Mux251~0_combout\) ) ) ) # ( \NxR.aluData2[0]~16_combout\ & ( !\Mux253~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & ((\Mux252~0_combout\))) # (\NxR.aluData2[1]~17_combout\ & 
-- (\Mux250~0_combout\)) ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( !\Mux253~0_combout\ & ( (\Mux251~0_combout\ & \NxR.aluData2[1]~17_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100010001000000111100111111011101110111010000001111001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux251~0_combout\,
	datab => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datac => \ALT_INV_Mux250~0_combout\,
	datad => \ALT_INV_Mux252~0_combout\,
	datae => \ALT_INV_NxR.aluData2[0]~16_combout\,
	dataf => \ALT_INV_Mux253~0_combout\,
	combout => \ShiftRight1~15_combout\);

-- Location: FF_X72_Y7_N7
\ShiftRight1~15_NEW_REG198\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~15_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~15_OTERM199\);

-- Location: MLABCELL_X78_Y9_N24
\ShiftRight1~19\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~19_combout\ = ( \ShiftRight1~17_OTERM267\ & ( \R.aluData2\(3) & ( (!\R.aluData2\(2)) # (\ShiftRight1~18_OTERM269\) ) ) ) # ( !\ShiftRight1~17_OTERM267\ & ( \R.aluData2\(3) & ( (\ShiftRight1~18_OTERM269\ & \R.aluData2\(2)) ) ) ) # ( 
-- \ShiftRight1~17_OTERM267\ & ( !\R.aluData2\(3) & ( (!\R.aluData2\(2) & ((\ShiftRight1~15_OTERM199\))) # (\R.aluData2\(2) & (\ShiftRight1~16_OTERM209\)) ) ) ) # ( !\ShiftRight1~17_OTERM267\ & ( !\R.aluData2\(3) & ( (!\R.aluData2\(2) & 
-- ((\ShiftRight1~15_OTERM199\))) # (\R.aluData2\(2) & (\ShiftRight1~16_OTERM209\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001111001111000000111100111100010001000100011101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~18_OTERM269\,
	datab => \ALT_INV_R.aluData2\(2),
	datac => \ALT_INV_ShiftRight1~16_OTERM209\,
	datad => \ALT_INV_ShiftRight1~15_OTERM199\,
	datae => \ALT_INV_ShiftRight1~17_OTERM267\,
	dataf => \ALT_INV_R.aluData2\(3),
	combout => \ShiftRight1~19_combout\);

-- Location: MLABCELL_X78_Y9_N42
\Selector31~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector31~1_combout\ = ( \R.aluOp.ALUOpSRA~q\ & ( \R.aluOp.ALUOpSRL~q\ & ( (!\R.aluData2\(4) & (((\ShiftRight1~19_combout\)))) # (\R.aluData2\(4) & (((\ShiftRight1~14_combout\)) # (\ShiftRight0~1_combout\))) ) ) ) # ( !\R.aluOp.ALUOpSRA~q\ & ( 
-- \R.aluOp.ALUOpSRL~q\ & ( (!\R.aluData2\(4) & ((\ShiftRight1~19_combout\))) # (\R.aluData2\(4) & (\ShiftRight0~1_combout\)) ) ) ) # ( \R.aluOp.ALUOpSRA~q\ & ( !\R.aluOp.ALUOpSRL~q\ & ( (!\R.aluData2\(4) & (\ShiftRight1~19_combout\)) # (\R.aluData2\(4) & 
-- ((\ShiftRight1~14_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000010100101111100011011000110110001101101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(4),
	datab => \ALT_INV_ShiftRight0~1_combout\,
	datac => \ALT_INV_ShiftRight1~19_combout\,
	datad => \ALT_INV_ShiftRight1~14_combout\,
	datae => \ALT_INV_R.aluOp.ALUOpSRA~q\,
	dataf => \ALT_INV_R.aluOp.ALUOpSRL~q\,
	combout => \Selector31~1_combout\);

-- Location: LABCELL_X83_Y5_N3
\Selector31~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector31~8_combout\ = ( \Selector31~4_combout\ & ( \Selector31~1_combout\ ) ) # ( !\Selector31~4_combout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111111111111111111100000000111111110000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \ALT_INV_Selector31~1_combout\,
	dataf => \ALT_INV_Selector31~4_combout\,
	combout => \Selector31~8_combout\);

-- Location: FF_X83_Y5_N4
\R.aluRes[1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector31~8_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(1));

-- Location: LABCELL_X81_Y9_N42
\vAluRes~1_RESYN1062\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~1_RESYN1062_BDD1063\ = ( \Selector31~1_combout\ & ( \Selector31~3_combout\ & ( (\R.aluRes\(1)) # (\R.aluCalc~q\) ) ) ) # ( !\Selector31~1_combout\ & ( \Selector31~3_combout\ & ( (!\R.aluCalc~q\ & \R.aluRes\(1)) ) ) ) # ( \Selector31~1_combout\ & 
-- ( !\Selector31~3_combout\ & ( (\R.aluRes\(1)) # (\R.aluCalc~q\) ) ) ) # ( !\Selector31~1_combout\ & ( !\Selector31~3_combout\ & ( (\R.aluRes\(1)) # (\R.aluCalc~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011111100111111001111110011111100001100000011000011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_R.aluRes\(1),
	datae => \ALT_INV_Selector31~1_combout\,
	dataf => \ALT_INV_Selector31~3_combout\,
	combout => \vAluRes~1_RESYN1062_BDD1063\);

-- Location: LABCELL_X81_Y9_N54
\vAluRes~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~1_combout\ = ( \Add2~5_sumout\ & ( \vAluRes~1_RESYN1062_BDD1063\ ) ) # ( !\Add2~5_sumout\ & ( \vAluRes~1_RESYN1062_BDD1063\ ) ) # ( \Add2~5_sumout\ & ( !\vAluRes~1_RESYN1062_BDD1063\ & ( (\R.aluCalc~q\ & (((\Add1~5_sumout\ & 
-- \R.aluOp.ALUOpAdd~q\)) # (\R.aluOp.ALUOpSub~q\))) ) ) ) # ( !\Add2~5_sumout\ & ( !\vAluRes~1_RESYN1062_BDD1063\ & ( (\Add1~5_sumout\ & (\R.aluCalc~q\ & \R.aluOp.ALUOpAdd~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000010001000000110001001111111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add1~5_sumout\,
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datad => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datae => \ALT_INV_Add2~5_sumout\,
	dataf => \ALT_INV_vAluRes~1_RESYN1062_BDD1063\,
	combout => \vAluRes~1_combout\);

-- Location: LABCELL_X83_Y5_N15
\Comb:vRegWriteData[1]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[1]~0_combout\ = ( \vAluRes~1_combout\ & ( (!\R.memToReg~q\) # ((\Mux222~0_combout\ & \avm_d_readdata[25]~input_o\)) ) ) # ( !\vAluRes~1_combout\ & ( (\R.memToReg~q\ & (\Mux222~0_combout\ & \avm_d_readdata[25]~input_o\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000100000001000000010000000110101011101010111010101110101011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.memToReg~q\,
	datab => \ALT_INV_Mux222~0_combout\,
	datac => \ALT_INV_avm_d_readdata[25]~input_o\,
	dataf => \ALT_INV_vAluRes~1_combout\,
	combout => \Comb:vRegWriteData[1]~0_combout\);

-- Location: FF_X83_Y5_N17
\R.regWriteData[1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vRegWriteData[1]~0_combout\,
	asdata => \R.curPC\(1),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(1));

-- Location: FF_X70_Y6_N38
\RegFile[15][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(1),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][1]~q\);

-- Location: LABCELL_X66_Y10_N27
\RegFile[14][1]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[14][1]~feeder_combout\ = ( \R.regWriteData\(1) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(1),
	combout => \RegFile[14][1]~feeder_combout\);

-- Location: FF_X66_Y10_N28
\RegFile[14][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[14][1]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][1]~q\);

-- Location: LABCELL_X63_Y8_N12
\RegFile[13][1]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[13][1]~feeder_combout\ = ( \R.regWriteData\(1) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(1),
	combout => \RegFile[13][1]~feeder_combout\);

-- Location: FF_X63_Y8_N13
\RegFile[13][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[13][1]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][1]~q\);

-- Location: FF_X63_Y8_N26
\RegFile[9][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(1),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][1]~q\);

-- Location: FF_X64_Y8_N49
\RegFile[10][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(1),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][1]~q\);

-- Location: FF_X70_Y6_N26
\RegFile[11][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(1),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][1]~q\);

-- Location: LABCELL_X63_Y8_N48
\RegFile[8][1]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[8][1]~feeder_combout\ = ( \R.regWriteData\(1) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(1),
	combout => \RegFile[8][1]~feeder_combout\);

-- Location: FF_X63_Y8_N49
\RegFile[8][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[8][1]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][1]~q\);

-- Location: LABCELL_X70_Y6_N24
\Mux121~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux121~14_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[8][1]~q\))) # (\R.curInst\(20) & (\RegFile[9][1]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & (\RegFile[10][1]~q\)) # (\R.curInst\(20) & ((\RegFile[11][1]~q\)))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001110111011101110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[9][1]~q\,
	datac => \ALT_INV_RegFile[10][1]~q\,
	datad => \ALT_INV_RegFile[11][1]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][1]~q\,
	combout => \Mux121~14_combout\);

-- Location: LABCELL_X66_Y7_N33
\RegFile[12][1]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[12][1]~feeder_combout\ = ( \R.regWriteData\(1) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(1),
	combout => \RegFile[12][1]~feeder_combout\);

-- Location: FF_X66_Y7_N34
\RegFile[12][1]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[12][1]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][1]~DUPLICATE_q\);

-- Location: LABCELL_X70_Y6_N36
\Mux121~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux121~1_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux121~14_combout\)))) # (\R.curInst\(22) & ((!\Mux121~14_combout\ & (\RegFile[12][1]~DUPLICATE_q\)) # (\Mux121~14_combout\ & ((\RegFile[13][1]~q\)))))) ) ) # ( \R.curInst\(21) & ( 
-- (!\R.curInst\(22) & ((((\Mux121~14_combout\))))) # (\R.curInst\(22) & (((!\Mux121~14_combout\ & ((\RegFile[14][1]~q\))) # (\Mux121~14_combout\ & (\RegFile[15][1]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111001100111111111101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][1]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[14][1]~q\,
	datad => \ALT_INV_RegFile[13][1]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux121~14_combout\,
	datag => \ALT_INV_RegFile[12][1]~DUPLICATE_q\,
	combout => \Mux121~1_combout\);

-- Location: FF_X70_Y4_N44
\RegFile[23][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(1),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][1]~q\);

-- Location: FF_X70_Y6_N32
\RegFile[21][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(1),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][1]~q\);

-- Location: FF_X75_Y8_N58
\RegFile[22][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(1),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][1]~q\);

-- Location: FF_X70_Y4_N20
\RegFile[19][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(1),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][1]~q\);

-- Location: FF_X70_Y4_N14
\RegFile[17][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(1),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][1]~q\);

-- Location: LABCELL_X71_Y4_N39
\RegFile[18][1]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[18][1]~feeder_combout\ = ( \R.regWriteData\(1) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(1),
	combout => \RegFile[18][1]~feeder_combout\);

-- Location: FF_X71_Y4_N40
\RegFile[18][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][1]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][1]~q\);

-- Location: FF_X75_Y4_N5
\RegFile[16][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(1),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][1]~q\);

-- Location: LABCELL_X70_Y4_N12
\Mux121~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux121~18_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[16][1]~q\))) # (\R.curInst\(20) & (\RegFile[17][1]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[18][1]~q\))) # (\R.curInst\(20) & (\RegFile[19][1]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[19][1]~q\,
	datab => \ALT_INV_RegFile[17][1]~q\,
	datac => \ALT_INV_RegFile[18][1]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][1]~q\,
	combout => \Mux121~18_combout\);

-- Location: FF_X77_Y8_N58
\RegFile[20][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(1),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][1]~q\);

-- Location: LABCELL_X70_Y6_N30
\Mux121~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux121~5_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux121~18_combout\)))) # (\R.curInst\(22) & ((!\Mux121~18_combout\ & ((\RegFile[20][1]~q\))) # (\Mux121~18_combout\ & (\RegFile[21][1]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux121~18_combout\)))) # (\R.curInst\(22) & ((!\Mux121~18_combout\ & ((\RegFile[22][1]~q\))) # (\Mux121~18_combout\ & (\RegFile[23][1]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[23][1]~q\,
	datab => \ALT_INV_RegFile[21][1]~q\,
	datac => \ALT_INV_RegFile[22][1]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux121~18_combout\,
	datag => \ALT_INV_RegFile[20][1]~q\,
	combout => \Mux121~5_combout\);

-- Location: FF_X66_Y6_N50
\RegFile[29][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(1),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][1]~q\);

-- Location: LABCELL_X68_Y8_N15
\RegFile[31][1]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[31][1]~feeder_combout\ = ( \R.regWriteData\(1) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(1),
	combout => \RegFile[31][1]~feeder_combout\);

-- Location: FF_X68_Y8_N16
\RegFile[31][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[31][1]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][1]~q\);

-- Location: FF_X66_Y6_N31
\RegFile[30][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(1),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][1]~q\);

-- Location: LABCELL_X67_Y4_N30
\RegFile[27][1]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[27][1]~feeder_combout\ = ( \R.regWriteData\(1) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(1),
	combout => \RegFile[27][1]~feeder_combout\);

-- Location: FF_X67_Y4_N31
\RegFile[27][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[27][1]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][1]~q\);

-- Location: LABCELL_X67_Y4_N3
\RegFile[26][1]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[26][1]~feeder_combout\ = ( \R.regWriteData\(1) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(1),
	combout => \RegFile[26][1]~feeder_combout\);

-- Location: FF_X67_Y4_N4
\RegFile[26][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[26][1]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][1]~q\);

-- Location: FF_X66_Y6_N8
\RegFile[25][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(1),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][1]~q\);

-- Location: LABCELL_X64_Y6_N12
\RegFile[24][1]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[24][1]~feeder_combout\ = ( \R.regWriteData\(1) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(1),
	combout => \RegFile[24][1]~feeder_combout\);

-- Location: FF_X64_Y6_N13
\RegFile[24][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[24][1]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][1]~q\);

-- Location: LABCELL_X66_Y6_N6
\Mux121~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux121~22_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & (\RegFile[24][1]~q\)) # (\R.curInst\(20) & ((\RegFile[25][1]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & ((\RegFile[26][1]~q\))) # (\R.curInst\(20) & (\RegFile[27][1]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110000110011111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[27][1]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[26][1]~q\,
	datad => \ALT_INV_RegFile[25][1]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][1]~q\,
	combout => \Mux121~22_combout\);

-- Location: LABCELL_X71_Y6_N18
\RegFile[28][1]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[28][1]~feeder_combout\ = ( \R.regWriteData\(1) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(1),
	combout => \RegFile[28][1]~feeder_combout\);

-- Location: FF_X71_Y6_N19
\RegFile[28][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[28][1]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][1]~q\);

-- Location: LABCELL_X66_Y6_N48
\Mux121~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux121~9_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux121~22_combout\)))) # (\R.curInst\(22) & ((!\Mux121~22_combout\ & ((\RegFile[28][1]~q\))) # (\Mux121~22_combout\ & (\RegFile[29][1]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux121~22_combout\)))) # (\R.curInst\(22) & ((!\Mux121~22_combout\ & ((\RegFile[30][1]~q\))) # (\Mux121~22_combout\ & (\RegFile[31][1]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[29][1]~q\,
	datab => \ALT_INV_RegFile[31][1]~q\,
	datac => \ALT_INV_RegFile[30][1]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux121~22_combout\,
	datag => \ALT_INV_RegFile[28][1]~q\,
	combout => \Mux121~9_combout\);

-- Location: FF_X67_Y7_N56
\RegFile[3][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(1),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][1]~q\);

-- Location: FF_X66_Y9_N37
\RegFile[2][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(1),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][1]~q\);

-- Location: FF_X66_Y9_N31
\RegFile[7][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(1),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][1]~q\);

-- Location: LABCELL_X63_Y7_N54
\RegFile[5][1]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[5][1]~feeder_combout\ = ( \R.regWriteData\(1) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(1),
	combout => \RegFile[5][1]~feeder_combout\);

-- Location: FF_X63_Y7_N55
\RegFile[5][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[5][1]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][1]~q\);

-- Location: FF_X67_Y5_N11
\RegFile[4][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(1),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][1]~q\);

-- Location: FF_X67_Y7_N49
\RegFile[6][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(1),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][1]~q\);

-- Location: LABCELL_X67_Y7_N48
\Mux121~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux121~0_combout\ = ( \RegFile[6][1]~q\ & ( \R.curInst\(21) & ( (!\R.curInst\(20)) # (\RegFile[7][1]~q\) ) ) ) # ( !\RegFile[6][1]~q\ & ( \R.curInst\(21) & ( (\RegFile[7][1]~q\ & \R.curInst\(20)) ) ) ) # ( \RegFile[6][1]~q\ & ( !\R.curInst\(21) & ( 
-- (!\R.curInst\(20) & ((\RegFile[4][1]~q\))) # (\R.curInst\(20) & (\RegFile[5][1]~q\)) ) ) ) # ( !\RegFile[6][1]~q\ & ( !\R.curInst\(21) & ( (!\R.curInst\(20) & ((\RegFile[4][1]~q\))) # (\R.curInst\(20) & (\RegFile[5][1]~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100110011000011110011001100000000010101011111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[7][1]~q\,
	datab => \ALT_INV_RegFile[5][1]~q\,
	datac => \ALT_INV_RegFile[4][1]~q\,
	datad => \ALT_INV_R.curInst\(20),
	datae => \ALT_INV_RegFile[6][1]~q\,
	dataf => \ALT_INV_R.curInst\(21),
	combout => \Mux121~0_combout\);

-- Location: LABCELL_X68_Y9_N42
\RegFile[1][1]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[1][1]~feeder_combout\ = ( \R.regWriteData\(1) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(1),
	combout => \RegFile[1][1]~feeder_combout\);

-- Location: FF_X68_Y9_N43
\RegFile[1][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[1][1]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][1]~q\);

-- Location: LABCELL_X67_Y7_N54
\Mux121~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux121~26_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (\RegFile[1][1]~q\ & (\R.curInst\(20)))) # (\R.curInst\(22) & (((\Mux121~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (((\RegFile[2][1]~q\)))) # 
-- (\R.curInst\(20) & (\RegFile[3][1]~q\)))) # (\R.curInst\(22) & ((((\Mux121~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001100000011000100010000110011001111110011111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][1]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[2][1]~q\,
	datad => \ALT_INV_R.curInst\(20),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux121~0_combout\,
	datag => \ALT_INV_RegFile[1][1]~q\,
	combout => \Mux121~26_combout\);

-- Location: LABCELL_X70_Y6_N6
\Mux121~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux121~13_combout\ = ( \Mux121~9_combout\ & ( \Mux121~26_combout\ & ( (!\R.curInst\(24) & ((!\R.curInst\(23)) # ((\Mux121~1_combout\)))) # (\R.curInst\(24) & (((\Mux121~5_combout\)) # (\R.curInst\(23)))) ) ) ) # ( !\Mux121~9_combout\ & ( 
-- \Mux121~26_combout\ & ( (!\R.curInst\(24) & ((!\R.curInst\(23)) # ((\Mux121~1_combout\)))) # (\R.curInst\(24) & (!\R.curInst\(23) & ((\Mux121~5_combout\)))) ) ) ) # ( \Mux121~9_combout\ & ( !\Mux121~26_combout\ & ( (!\R.curInst\(24) & (\R.curInst\(23) & 
-- (\Mux121~1_combout\))) # (\R.curInst\(24) & (((\Mux121~5_combout\)) # (\R.curInst\(23)))) ) ) ) # ( !\Mux121~9_combout\ & ( !\Mux121~26_combout\ & ( (!\R.curInst\(24) & (\R.curInst\(23) & (\Mux121~1_combout\))) # (\R.curInst\(24) & (!\R.curInst\(23) & 
-- ((\Mux121~5_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001001000110000100110101011110001010110011101001101111011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(24),
	datab => \ALT_INV_R.curInst\(23),
	datac => \ALT_INV_Mux121~1_combout\,
	datad => \ALT_INV_Mux121~5_combout\,
	datae => \ALT_INV_Mux121~9_combout\,
	dataf => \ALT_INV_Mux121~26_combout\,
	combout => \Mux121~13_combout\);

-- Location: LABCELL_X74_Y6_N6
\NxR.aluData2[1]~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[1]~17_combout\ = ( \Mux121~13_combout\ & ( (!\vAluSrc2~1_combout\) # ((\Equal4~1_combout\ & \Mux153~0_combout\)) ) ) # ( !\Mux121~13_combout\ & ( (\Equal4~1_combout\ & (\Mux153~0_combout\ & \vAluSrc2~1_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000011000000000000001111111111000000111111111100000011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Equal4~1_combout\,
	datac => \ALT_INV_Mux153~0_combout\,
	datad => \ALT_INV_vAluSrc2~1_combout\,
	dataf => \ALT_INV_Mux121~13_combout\,
	combout => \NxR.aluData2[1]~17_combout\);

-- Location: FF_X75_Y6_N40
\R.aluData2[1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \NxR.aluData2[1]~17_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData2\(1));

-- Location: LABCELL_X77_Y9_N12
\Selector18~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector18~0_combout\ = ( \R.aluData1\(30) & ( \R.aluData1\(31) & ( ((\R.aluOp.ALUOpSRL~q\ & !\R.aluData2\(1))) # (\R.aluOp.ALUOpSRA~q\) ) ) ) # ( !\R.aluData1\(30) & ( \R.aluData1\(31) & ( (!\R.aluData2\(1) & (\R.aluData2\(0) & ((\R.aluOp.ALUOpSRA~q\) # 
-- (\R.aluOp.ALUOpSRL~q\)))) # (\R.aluData2\(1) & (((\R.aluOp.ALUOpSRA~q\)))) ) ) ) # ( \R.aluData1\(30) & ( !\R.aluData1\(31) & ( (!\R.aluData2\(0) & (!\R.aluData2\(1) & ((\R.aluOp.ALUOpSRA~q\) # (\R.aluOp.ALUOpSRL~q\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000001000001010000000010000010111110011000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(0),
	datab => \ALT_INV_R.aluOp.ALUOpSRL~q\,
	datac => \ALT_INV_R.aluData2\(1),
	datad => \ALT_INV_R.aluOp.ALUOpSRA~q\,
	datae => \ALT_INV_R.aluData1\(30),
	dataf => \ALT_INV_R.aluData1\(31),
	combout => \Selector18~0_combout\);

-- Location: LABCELL_X74_Y9_N27
\Selector18~1_RTM0433\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector18~1_RTM0433_combout\ = ( \Mux240~0_combout\ & ( \R.aluOp.ALUOpAnd_OTERM357\ & ( ((\NxR.aluData2[14]~7_combout\) # (\R.aluOp.ALUOpXor_OTERM355\)) # (\R.aluOp.ALUOpOr_OTERM353\) ) ) ) # ( !\Mux240~0_combout\ & ( \R.aluOp.ALUOpAnd_OTERM357\ & ( 
-- (\NxR.aluData2[14]~7_combout\ & ((\R.aluOp.ALUOpXor_OTERM355\) # (\R.aluOp.ALUOpOr_OTERM353\))) ) ) ) # ( \Mux240~0_combout\ & ( !\R.aluOp.ALUOpAnd_OTERM357\ & ( ((\R.aluOp.ALUOpXor_OTERM355\ & !\NxR.aluData2[14]~7_combout\)) # 
-- (\R.aluOp.ALUOpOr_OTERM353\) ) ) ) # ( !\Mux240~0_combout\ & ( !\R.aluOp.ALUOpAnd_OTERM357\ & ( (\NxR.aluData2[14]~7_combout\ & ((\R.aluOp.ALUOpXor_OTERM355\) # (\R.aluOp.ALUOpOr_OTERM353\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001011111010111110101010100000000010111110101111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpOr_OTERM353\,
	datac => \ALT_INV_R.aluOp.ALUOpXor_OTERM355\,
	datad => \ALT_INV_NxR.aluData2[14]~7_combout\,
	datae => \ALT_INV_Mux240~0_combout\,
	dataf => \ALT_INV_R.aluOp.ALUOpAnd_OTERM357\,
	combout => \Selector18~1_RTM0433_combout\);

-- Location: FF_X74_Y9_N28
\Selector18~1_NEW_REG430\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector18~1_RTM0433_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector18~1_OTERM431\);

-- Location: LABCELL_X77_Y9_N42
\Selector18~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector18~2_combout\ = ( \Selector20~0_OTERM769\ & ( (!\R.aluData2\(4) & !\Selector18~1_OTERM431\) ) ) # ( !\Selector20~0_OTERM769\ & ( (!\Selector18~1_OTERM431\ & ((!\R.aluData2\(4)) # ((!\Selector18~0_combout\) # 
-- (\ShiftRight0~7_OTERM233DUPLICATE_q\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1110111100000000111011110000000010101010000000001010101000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(4),
	datab => \ALT_INV_Selector18~0_combout\,
	datac => \ALT_INV_ShiftRight0~7_OTERM233DUPLICATE_q\,
	datad => \ALT_INV_Selector18~1_OTERM431\,
	dataf => \ALT_INV_Selector20~0_OTERM769\,
	combout => \Selector18~2_combout\);

-- Location: MLABCELL_X78_Y7_N6
\ShiftLeft0~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~21_combout\ = ( \ShiftLeft0~20_OTERM291\ & ( \R.aluData2\(3) & ( (!\R.aluData2\(2) & ((\ShiftLeft0~8_OTERM207\))) # (\R.aluData2\(2) & (\ShiftLeft0~2_OTERM221\)) ) ) ) # ( !\ShiftLeft0~20_OTERM291\ & ( \R.aluData2\(3) & ( (!\R.aluData2\(2) & 
-- ((\ShiftLeft0~8_OTERM207\))) # (\R.aluData2\(2) & (\ShiftLeft0~2_OTERM221\)) ) ) ) # ( \ShiftLeft0~20_OTERM291\ & ( !\R.aluData2\(3) & ( (!\R.aluData2\(2)) # (\ShiftLeft0~13_OTERM285\) ) ) ) # ( !\ShiftLeft0~20_OTERM291\ & ( !\R.aluData2\(3) & ( 
-- (\ShiftLeft0~13_OTERM285\ & \R.aluData2\(2)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100010001110111011101110100000011110011110000001111001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~13_OTERM285\,
	datab => \ALT_INV_R.aluData2\(2),
	datac => \ALT_INV_ShiftLeft0~2_OTERM221\,
	datad => \ALT_INV_ShiftLeft0~8_OTERM207\,
	datae => \ALT_INV_ShiftLeft0~20_OTERM291\,
	dataf => \ALT_INV_R.aluData2\(3),
	combout => \ShiftLeft0~21_combout\);

-- Location: MLABCELL_X82_Y6_N36
\ShiftRight1~53\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~53_combout\ = ( \R.aluData2\(2) & ( \ShiftRight1~27_OTERM19\ & ( (\ShiftRight1~25_OTERM277\) # (\R.aluData2\(3)) ) ) ) # ( !\R.aluData2\(2) & ( \ShiftRight1~27_OTERM19\ & ( (!\R.aluData2\(3) & ((\ShiftRight1~23_OTERM275\))) # (\R.aluData2\(3) 
-- & (\ShiftRight1~26_OTERM37\)) ) ) ) # ( \R.aluData2\(2) & ( !\ShiftRight1~27_OTERM19\ & ( (!\R.aluData2\(3) & \ShiftRight1~25_OTERM277\) ) ) ) # ( !\R.aluData2\(2) & ( !\ShiftRight1~27_OTERM19\ & ( (!\R.aluData2\(3) & ((\ShiftRight1~23_OTERM275\))) # 
-- (\R.aluData2\(3) & (\ShiftRight1~26_OTERM37\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010110101111001000100010001000000101101011110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(3),
	datab => \ALT_INV_ShiftRight1~25_OTERM277\,
	datac => \ALT_INV_ShiftRight1~26_OTERM37\,
	datad => \ALT_INV_ShiftRight1~23_OTERM275\,
	datae => \ALT_INV_R.aluData2\(2),
	dataf => \ALT_INV_ShiftRight1~27_OTERM19\,
	combout => \ShiftRight1~53_combout\);

-- Location: LABCELL_X83_Y7_N57
\Selector18~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector18~3_combout\ = ( \Selector27~0_OTERM385\ & ( \ShiftRight1~53_combout\ & ( (!\Selector31~5_OTERM599\ & (\Selector18~2_combout\ & !\ShiftLeft0~21_combout\)) ) ) ) # ( !\Selector27~0_OTERM385\ & ( \ShiftRight1~53_combout\ & ( 
-- (!\Selector31~5_OTERM599\ & \Selector18~2_combout\) ) ) ) # ( \Selector27~0_OTERM385\ & ( !\ShiftRight1~53_combout\ & ( (\Selector18~2_combout\ & !\ShiftLeft0~21_combout\) ) ) ) # ( !\Selector27~0_OTERM385\ & ( !\ShiftRight1~53_combout\ & ( 
-- \Selector18~2_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110011001100000011000000100010001000100010000000100000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector31~5_OTERM599\,
	datab => \ALT_INV_Selector18~2_combout\,
	datac => \ALT_INV_ShiftLeft0~21_combout\,
	datae => \ALT_INV_Selector27~0_OTERM385\,
	dataf => \ALT_INV_ShiftRight1~53_combout\,
	combout => \Selector18~3_combout\);

-- Location: MLABCELL_X78_Y3_N45
\Selector18~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector18~4_combout\ = ( \Add2~57_sumout\ & ( ((\R.aluOp.ALUOpAdd~q\ & \Add1~57_sumout\)) # (\R.aluOp.ALUOpSub~q\) ) ) # ( !\Add2~57_sumout\ & ( (\R.aluOp.ALUOpAdd~q\ & \Add1~57_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101000001010000010100000101111111110000010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datac => \ALT_INV_Add1~57_sumout\,
	datad => \ALT_INV_R.aluOp.ALUOpSub~q\,
	dataf => \ALT_INV_Add2~57_sumout\,
	combout => \Selector18~4_combout\);

-- Location: MLABCELL_X78_Y3_N36
\Comb:vJumpAdr[14]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[14]~0_combout\ = ( \R.aluCalc~q\ & ( \Add3~57_sumout\ & ( (!\Selector18~3_combout\) # ((!\Equal4~2_combout\) # (\Selector18~4_combout\)) ) ) ) # ( !\R.aluCalc~q\ & ( \Add3~57_sumout\ & ( (!\Equal4~2_combout\) # (\R.aluRes\(14)) ) ) ) # ( 
-- \R.aluCalc~q\ & ( !\Add3~57_sumout\ & ( (\Equal4~2_combout\ & ((!\Selector18~3_combout\) # (\Selector18~4_combout\))) ) ) ) # ( !\R.aluCalc~q\ & ( !\Add3~57_sumout\ & ( (\Equal4~2_combout\ & \R.aluRes\(14)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011001000100011001111001111110011111110111011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector18~3_combout\,
	datab => \ALT_INV_Equal4~2_combout\,
	datac => \ALT_INV_R.aluRes\(14),
	datad => \ALT_INV_Selector18~4_combout\,
	datae => \ALT_INV_R.aluCalc~q\,
	dataf => \ALT_INV_Add3~57_sumout\,
	combout => \Comb:vJumpAdr[14]~0_combout\);

-- Location: FF_X78_Y3_N37
\R.curPC[14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[14]~0_combout\,
	asdata => \Add0~49_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(14));

-- Location: LABCELL_X63_Y6_N30
\Mux76~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux76~14_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[8][14]~q\))) # (\R.curInst\(15) & (\RegFile[9][14]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & (\RegFile[10][14]~q\)) # (\R.curInst\(15) & ((\RegFile[11][14]~q\)))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001110111011101110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[9][14]~q\,
	datac => \ALT_INV_RegFile[10][14]~q\,
	datad => \ALT_INV_RegFile[11][14]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][14]~q\,
	combout => \Mux76~14_combout\);

-- Location: LABCELL_X63_Y6_N48
\Mux76~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux76~1_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux76~14_combout\)))) # (\R.curInst\(17) & ((!\Mux76~14_combout\ & (\RegFile[12][14]~q\)) # (\Mux76~14_combout\ & ((\RegFile[13][14]~q\)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) 
-- & ((((\Mux76~14_combout\))))) # (\R.curInst\(17) & (((!\Mux76~14_combout\ & ((\RegFile[14][14]~q\))) # (\Mux76~14_combout\ & (\RegFile[15][14]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111001100111111111101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][14]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[14][14]~q\,
	datad => \ALT_INV_RegFile[13][14]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux76~14_combout\,
	datag => \ALT_INV_RegFile[12][14]~q\,
	combout => \Mux76~1_combout\);

-- Location: LABCELL_X63_Y6_N24
\Mux76~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux76~22_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[24][14]~q\))) # (\R.curInst\(15) & (\RegFile[25][14]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[26][14]~q\))) # (\R.curInst\(15) & (\RegFile[27][14]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[27][14]~q\,
	datab => \ALT_INV_RegFile[25][14]~q\,
	datac => \ALT_INV_RegFile[26][14]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][14]~q\,
	combout => \Mux76~22_combout\);

-- Location: LABCELL_X63_Y6_N6
\Mux76~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux76~9_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux76~22_combout\)))) # (\R.curInst\(17) & ((!\Mux76~22_combout\ & ((\RegFile[28][14]~q\))) # (\Mux76~22_combout\ & (\RegFile[29][14]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux76~22_combout\)))) # (\R.curInst\(17) & ((!\Mux76~22_combout\ & ((\RegFile[30][14]~q\))) # (\Mux76~22_combout\ & (\RegFile[31][14]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[29][14]~q\,
	datab => \ALT_INV_RegFile[31][14]~q\,
	datac => \ALT_INV_RegFile[30][14]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux76~22_combout\,
	datag => \ALT_INV_RegFile[28][14]~q\,
	combout => \Mux76~9_combout\);

-- Location: LABCELL_X64_Y2_N42
\Mux76~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux76~18_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[16][14]~q\))) # (\R.curInst\(15) & (\RegFile[17][14]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[18][14]~q\))) # (\R.curInst\(15) & (\RegFile[19][14]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[19][14]~q\,
	datab => \ALT_INV_RegFile[17][14]~q\,
	datac => \ALT_INV_RegFile[18][14]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][14]~q\,
	combout => \Mux76~18_combout\);

-- Location: LABCELL_X64_Y2_N36
\Mux76~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux76~5_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux76~18_combout\)))) # (\R.curInst\(17) & ((!\Mux76~18_combout\ & (\RegFile[20][14]~q\)) # (\Mux76~18_combout\ & ((\RegFile[21][14]~q\)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) 
-- & ((((\Mux76~18_combout\))))) # (\R.curInst\(17) & (((!\Mux76~18_combout\ & ((\RegFile[22][14]~q\))) # (\Mux76~18_combout\ & (\RegFile[23][14]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111001100111111111101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[23][14]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[22][14]~q\,
	datad => \ALT_INV_RegFile[21][14]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux76~18_combout\,
	datag => \ALT_INV_RegFile[20][14]~q\,
	combout => \Mux76~5_combout\);

-- Location: LABCELL_X62_Y8_N12
\Mux76~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux76~0_combout\ = ( \RegFile[7][14]~q\ & ( \R.curInst\(16) & ( (\R.curInst\(15)) # (\RegFile[6][14]~q\) ) ) ) # ( !\RegFile[7][14]~q\ & ( \R.curInst\(16) & ( (\RegFile[6][14]~q\ & !\R.curInst\(15)) ) ) ) # ( \RegFile[7][14]~q\ & ( !\R.curInst\(16) & ( 
-- (!\R.curInst\(15) & ((\RegFile[4][14]~q\))) # (\R.curInst\(15) & (\RegFile[5][14]~q\)) ) ) ) # ( !\RegFile[7][14]~q\ & ( !\R.curInst\(16) & ( (!\R.curInst\(15) & ((\RegFile[4][14]~q\))) # (\R.curInst\(15) & (\RegFile[5][14]~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100110011000011110011001101010101000000000101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[6][14]~q\,
	datab => \ALT_INV_RegFile[5][14]~q\,
	datac => \ALT_INV_RegFile[4][14]~q\,
	datad => \ALT_INV_R.curInst\(15),
	datae => \ALT_INV_RegFile[7][14]~q\,
	dataf => \ALT_INV_R.curInst\(16),
	combout => \Mux76~0_combout\);

-- Location: FF_X59_Y7_N58
\RegFile[1][14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[1][14]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][14]~q\);

-- Location: LABCELL_X62_Y8_N30
\Mux76~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux76~26_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (\R.curInst\(15) & (\RegFile[1][14]~q\))) # (\R.curInst\(17) & (((\Mux76~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & ((!\R.curInst\(15) & (((\RegFile[2][14]~q\)))) # 
-- (\R.curInst\(15) & (\RegFile[3][14]~q\)))) # (\R.curInst\(17) & ((((\Mux76~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000000000110110000000000000101111111110001101111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(15),
	datab => \ALT_INV_RegFile[3][14]~q\,
	datac => \ALT_INV_RegFile[2][14]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux76~0_combout\,
	datag => \ALT_INV_RegFile[1][14]~q\,
	combout => \Mux76~26_combout\);

-- Location: LABCELL_X63_Y6_N36
\Mux76~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux76~13_combout\ = ( \Mux76~5_combout\ & ( \Mux76~26_combout\ & ( (!\R.curInst\(18)) # ((!\R.curInst\(19) & (\Mux76~1_combout\)) # (\R.curInst\(19) & ((\Mux76~9_combout\)))) ) ) ) # ( !\Mux76~5_combout\ & ( \Mux76~26_combout\ & ( (!\R.curInst\(18) & 
-- (!\R.curInst\(19))) # (\R.curInst\(18) & ((!\R.curInst\(19) & (\Mux76~1_combout\)) # (\R.curInst\(19) & ((\Mux76~9_combout\))))) ) ) ) # ( \Mux76~5_combout\ & ( !\Mux76~26_combout\ & ( (!\R.curInst\(18) & (\R.curInst\(19))) # (\R.curInst\(18) & 
-- ((!\R.curInst\(19) & (\Mux76~1_combout\)) # (\R.curInst\(19) & ((\Mux76~9_combout\))))) ) ) ) # ( !\Mux76~5_combout\ & ( !\Mux76~26_combout\ & ( (\R.curInst\(18) & ((!\R.curInst\(19) & (\Mux76~1_combout\)) # (\R.curInst\(19) & ((\Mux76~9_combout\))))) ) ) 
-- )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010000010101001001100011011110001100100111011010111010111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(18),
	datab => \ALT_INV_R.curInst\(19),
	datac => \ALT_INV_Mux76~1_combout\,
	datad => \ALT_INV_Mux76~9_combout\,
	datae => \ALT_INV_Mux76~5_combout\,
	dataf => \ALT_INV_Mux76~26_combout\,
	combout => \Mux76~13_combout\);

-- Location: LABCELL_X73_Y6_N36
\Mux240~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux240~0_combout\ = ( \Mux76~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC\(14)))) ) ) # ( !\Mux76~13_combout\ & ( (\R.curPC\(14) & (\vAluSrc1~2_combout\ & !\vAluSrc1~1_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000000000000110000000011110011000000001111001100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.curPC\(14),
	datac => \ALT_INV_vAluSrc1~2_combout\,
	datad => \ALT_INV_vAluSrc1~1_combout\,
	dataf => \ALT_INV_Mux76~13_combout\,
	combout => \Mux240~0_combout\);

-- Location: LABCELL_X73_Y6_N6
\ShiftLeft0~24\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~24_combout\ = ( \Mux239~0_combout\ & ( \Mux238~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\) # ((!\NxR.aluData2[0]~16_combout\ & (\Mux240~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & ((\Mux241~0_combout\)))) ) ) ) # ( !\Mux239~0_combout\ & 
-- ( \Mux238~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (((!\NxR.aluData2[1]~17_combout\)) # (\Mux240~0_combout\))) # (\NxR.aluData2[0]~16_combout\ & (((\NxR.aluData2[1]~17_combout\ & \Mux241~0_combout\)))) ) ) ) # ( \Mux239~0_combout\ & ( 
-- !\Mux238~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (\Mux240~0_combout\ & (\NxR.aluData2[1]~17_combout\))) # (\NxR.aluData2[0]~16_combout\ & (((!\NxR.aluData2[1]~17_combout\) # (\Mux241~0_combout\)))) ) ) ) # ( !\Mux239~0_combout\ & ( 
-- !\Mux238~0_combout\ & ( (\NxR.aluData2[1]~17_combout\ & ((!\NxR.aluData2[0]~16_combout\ & (\Mux240~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & ((\Mux241~0_combout\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001000000111010100100101011110100010101001111111001011110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datab => \ALT_INV_Mux240~0_combout\,
	datac => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datad => \ALT_INV_Mux241~0_combout\,
	datae => \ALT_INV_Mux239~0_combout\,
	dataf => \ALT_INV_Mux238~0_combout\,
	combout => \ShiftLeft0~24_combout\);

-- Location: FF_X73_Y6_N7
\ShiftLeft0~24_NEW_REG292\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~24_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~24_OTERM293\);

-- Location: LABCELL_X81_Y8_N42
\ShiftLeft0~33\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~33_combout\ = ( \ShiftLeft0~10_OTERM211\ & ( \ShiftLeft0~32_OTERM297\ & ( (!\R.aluData2\(3) & (((!\R.aluData2\(2))) # (\ShiftLeft0~24_OTERM293\))) # (\R.aluData2\(3) & (((\ShiftLeft0~16_OTERM287\) # (\R.aluData2\(2))))) ) ) ) # ( 
-- !\ShiftLeft0~10_OTERM211\ & ( \ShiftLeft0~32_OTERM297\ & ( (!\R.aluData2\(3) & (((!\R.aluData2\(2))) # (\ShiftLeft0~24_OTERM293\))) # (\R.aluData2\(3) & (((!\R.aluData2\(2) & \ShiftLeft0~16_OTERM287\)))) ) ) ) # ( \ShiftLeft0~10_OTERM211\ & ( 
-- !\ShiftLeft0~32_OTERM297\ & ( (!\R.aluData2\(3) & (\ShiftLeft0~24_OTERM293\ & (\R.aluData2\(2)))) # (\R.aluData2\(3) & (((\ShiftLeft0~16_OTERM287\) # (\R.aluData2\(2))))) ) ) ) # ( !\ShiftLeft0~10_OTERM211\ & ( !\ShiftLeft0~32_OTERM297\ & ( 
-- (!\R.aluData2\(3) & (\ShiftLeft0~24_OTERM293\ & (\R.aluData2\(2)))) # (\R.aluData2\(3) & (((!\R.aluData2\(2) & \ShiftLeft0~16_OTERM287\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010000110100000001110011011111000100111101001100011111110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~24_OTERM293\,
	datab => \ALT_INV_R.aluData2\(3),
	datac => \ALT_INV_R.aluData2\(2),
	datad => \ALT_INV_ShiftLeft0~16_OTERM287\,
	datae => \ALT_INV_ShiftLeft0~10_OTERM211\,
	dataf => \ALT_INV_ShiftLeft0~32_OTERM297\,
	combout => \ShiftLeft0~33_combout\);

-- Location: LABCELL_X81_Y8_N12
\Selector12~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector12~0_combout\ = ( \ShiftRight1~3_OTERM13\ & ( \R.aluData2\(2) & ( (\ShiftRight1~2_OTERM49\ & (!\R.aluData2\(3) & \R.aluOp.ALUOpSRL~q\)) ) ) ) # ( !\ShiftRight1~3_OTERM13\ & ( \R.aluData2\(2) & ( (\ShiftRight1~2_OTERM49\ & (!\R.aluData2\(3) & 
-- \R.aluOp.ALUOpSRL~q\)) ) ) ) # ( \ShiftRight1~3_OTERM13\ & ( !\R.aluData2\(2) & ( (\R.aluOp.ALUOpSRL~q\ & ((\ShiftRight1~1_OTERM33\) # (\R.aluData2\(3)))) ) ) ) # ( !\ShiftRight1~3_OTERM13\ & ( !\R.aluData2\(2) & ( (!\R.aluData2\(3) & 
-- (\R.aluOp.ALUOpSRL~q\ & \ShiftRight1~1_OTERM33\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000001100000000110000111100000100000001000000010000000100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~2_OTERM49\,
	datab => \ALT_INV_R.aluData2\(3),
	datac => \ALT_INV_R.aluOp.ALUOpSRL~q\,
	datad => \ALT_INV_ShiftRight1~1_OTERM33\,
	datae => \ALT_INV_ShiftRight1~3_OTERM13\,
	dataf => \ALT_INV_R.aluData2\(2),
	combout => \Selector12~0_combout\);

-- Location: LABCELL_X75_Y8_N15
\ShiftRight1~39\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~39_combout\ = ( \R.aluData1\(31) & ( \R.aluData2\(2) & ( (\ShiftRight1~2_OTERM49\) # (\R.aluData2\(3)) ) ) ) # ( !\R.aluData1\(31) & ( \R.aluData2\(2) & ( (!\R.aluData2\(3) & \ShiftRight1~2_OTERM49\) ) ) ) # ( \R.aluData1\(31) & ( 
-- !\R.aluData2\(2) & ( (!\R.aluData2\(3) & ((\ShiftRight1~1_OTERM33\))) # (\R.aluData2\(3) & (\ShiftRight1~3_OTERM13\)) ) ) ) # ( !\R.aluData1\(31) & ( !\R.aluData2\(2) & ( (!\R.aluData2\(3) & ((\ShiftRight1~1_OTERM33\))) # (\R.aluData2\(3) & 
-- (\ShiftRight1~3_OTERM13\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000111011101000100011101110100001100000011000011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~3_OTERM13\,
	datab => \ALT_INV_R.aluData2\(3),
	datac => \ALT_INV_ShiftRight1~2_OTERM49\,
	datad => \ALT_INV_ShiftRight1~1_OTERM33\,
	datae => \ALT_INV_R.aluData1\(31),
	dataf => \ALT_INV_R.aluData2\(2),
	combout => \ShiftRight1~39_combout\);

-- Location: MLABCELL_X82_Y8_N57
\Selector12~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector12~1_combout\ = ( \Selector12~0_combout\ & ( \ShiftRight1~39_combout\ & ( !\R.aluData2\(4) ) ) ) # ( !\Selector12~0_combout\ & ( \ShiftRight1~39_combout\ & ( (!\R.aluData2\(4) & (((\R.aluOp.ALUOpSLL~q\ & \ShiftLeft0~33_combout\)) # 
-- (\R.aluOp.ALUOpSRA~q\))) ) ) ) # ( \Selector12~0_combout\ & ( !\ShiftRight1~39_combout\ & ( !\R.aluData2\(4) ) ) ) # ( !\Selector12~0_combout\ & ( !\ShiftRight1~39_combout\ & ( (\R.aluOp.ALUOpSLL~q\ & (\ShiftLeft0~33_combout\ & !\R.aluData2\(4))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000000010000111100001111000000010000111100001111000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpSLL~q\,
	datab => \ALT_INV_ShiftLeft0~33_combout\,
	datac => \ALT_INV_R.aluData2\(4),
	datad => \ALT_INV_R.aluOp.ALUOpSRA~q\,
	datae => \ALT_INV_Selector12~0_combout\,
	dataf => \ALT_INV_ShiftRight1~39_combout\,
	combout => \Selector12~1_combout\);

-- Location: MLABCELL_X78_Y8_N24
\Selector12~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector12~5_combout\ = ( \Selector12~4_combout\ & ( \Add2~81_sumout\ & ( (((\R.aluOp.ALUOpAdd~q\ & \Add1~81_sumout\)) # (\R.aluOp.ALUOpSub~q\)) # (\Selector12~1_combout\) ) ) ) # ( !\Selector12~4_combout\ & ( \Add2~81_sumout\ ) ) # ( 
-- \Selector12~4_combout\ & ( !\Add2~81_sumout\ & ( ((\R.aluOp.ALUOpAdd~q\ & \Add1~81_sumout\)) # (\Selector12~1_combout\) ) ) ) # ( !\Selector12~4_combout\ & ( !\Add2~81_sumout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111010101010111011111111111111111110101111101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector12~1_combout\,
	datab => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datac => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datad => \ALT_INV_Add1~81_sumout\,
	datae => \ALT_INV_Selector12~4_combout\,
	dataf => \ALT_INV_Add2~81_sumout\,
	combout => \Selector12~5_combout\);

-- Location: FF_X78_Y8_N26
\R.aluRes[20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector12~5_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(20));

-- Location: MLABCELL_X78_Y8_N0
\Comb:vJumpAdr[20]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[20]~0_combout\ = ( \Add3~81_sumout\ & ( (!\Equal4~2_combout\) # ((!\R.aluCalc~q\ & (\R.aluRes\(20))) # (\R.aluCalc~q\ & ((\Selector12~5_combout\)))) ) ) # ( !\Add3~81_sumout\ & ( (\Equal4~2_combout\ & ((!\R.aluCalc~q\ & (\R.aluRes\(20))) # 
-- (\R.aluCalc~q\ & ((\Selector12~5_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001000111000000000100011111111111010001111111111101000111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluRes\(20),
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_Selector12~5_combout\,
	datad => \ALT_INV_Equal4~2_combout\,
	dataf => \ALT_INV_Add3~81_sumout\,
	combout => \Comb:vJumpAdr[20]~0_combout\);

-- Location: FF_X78_Y8_N1
\R.curPC[20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[20]~0_combout\,
	asdata => \Add0~73_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(20));

-- Location: LABCELL_X68_Y3_N30
\Mux70~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux70~0_combout\ = ( \RegFile[7][20]~q\ & ( \R.curInst\(15) & ( (\RegFile[5][20]~q\) # (\R.curInst\(16)) ) ) ) # ( !\RegFile[7][20]~q\ & ( \R.curInst\(15) & ( (!\R.curInst\(16) & \RegFile[5][20]~q\) ) ) ) # ( \RegFile[7][20]~q\ & ( !\R.curInst\(15) & ( 
-- (!\R.curInst\(16) & ((\RegFile[4][20]~q\))) # (\R.curInst\(16) & (\RegFile[6][20]~q\)) ) ) ) # ( !\RegFile[7][20]~q\ & ( !\R.curInst\(15) & ( (!\R.curInst\(16) & ((\RegFile[4][20]~q\))) # (\R.curInst\(16) & (\RegFile[6][20]~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001110100011101000111010001110100000000110011000011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[6][20]~q\,
	datab => \ALT_INV_R.curInst\(16),
	datac => \ALT_INV_RegFile[4][20]~q\,
	datad => \ALT_INV_RegFile[5][20]~q\,
	datae => \ALT_INV_RegFile[7][20]~q\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux70~0_combout\);

-- Location: FF_X72_Y3_N55
\RegFile[1][20]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[1][20]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][20]~DUPLICATE_q\);

-- Location: LABCELL_X67_Y3_N12
\Mux70~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux70~26_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (\R.curInst\(15) & (\RegFile[1][20]~DUPLICATE_q\))) # (\R.curInst\(17) & (((\Mux70~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & ((!\R.curInst\(15) & 
-- (((\RegFile[2][20]~q\)))) # (\R.curInst\(15) & (\RegFile[3][20]~q\)))) # (\R.curInst\(17) & ((((\Mux70~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000000000111010000000000000011111111110001110111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][20]~q\,
	datab => \ALT_INV_R.curInst\(15),
	datac => \ALT_INV_RegFile[2][20]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux70~0_combout\,
	datag => \ALT_INV_RegFile[1][20]~DUPLICATE_q\,
	combout => \Mux70~26_combout\);

-- Location: FF_X63_Y3_N50
\RegFile[14][20]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(20),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][20]~q\);

-- Location: LABCELL_X63_Y1_N36
\Mux70~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux70~14_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[8][20]~q\))) # (\R.curInst\(15) & (\RegFile[9][20]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[10][20]~q\))) # (\R.curInst\(15) & (\RegFile[11][20]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[11][20]~q\,
	datab => \ALT_INV_RegFile[9][20]~q\,
	datac => \ALT_INV_RegFile[10][20]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][20]~q\,
	combout => \Mux70~14_combout\);

-- Location: LABCELL_X63_Y3_N24
\Mux70~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux70~1_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux70~14_combout\)))) # (\R.curInst\(17) & ((!\Mux70~14_combout\ & (\RegFile[12][20]~q\)) # (\Mux70~14_combout\ & ((\RegFile[13][20]~q\)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) 
-- & ((((\Mux70~14_combout\))))) # (\R.curInst\(17) & (((!\Mux70~14_combout\ & ((\RegFile[14][20]~q\))) # (\Mux70~14_combout\ & (\RegFile[15][20]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111001100111111111101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][20]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[14][20]~q\,
	datad => \ALT_INV_RegFile[13][20]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux70~14_combout\,
	datag => \ALT_INV_RegFile[12][20]~q\,
	combout => \Mux70~1_combout\);

-- Location: LABCELL_X66_Y2_N30
\Mux70~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux70~22_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[24][20]~q\))) # (\R.curInst\(15) & (\RegFile[25][20]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & (\RegFile[26][20]~q\)) # (\R.curInst\(15) & ((\RegFile[27][20]~q\))))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[25][20]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[26][20]~q\,
	datad => \ALT_INV_RegFile[27][20]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][20]~q\,
	combout => \Mux70~22_combout\);

-- Location: LABCELL_X66_Y3_N6
\Mux70~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux70~9_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux70~22_combout\))))) # (\R.curInst\(17) & (((!\Mux70~22_combout\ & (\RegFile[28][20]~q\)) # (\Mux70~22_combout\ & ((\RegFile[29][20]~q\)))))) ) ) # ( \R.curInst\(16) & ( 
-- (!\R.curInst\(17) & ((((\Mux70~22_combout\))))) # (\R.curInst\(17) & (((!\Mux70~22_combout\ & ((\RegFile[30][20]~q\))) # (\Mux70~22_combout\ & (\RegFile[31][20]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110101010111111111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[31][20]~q\,
	datac => \ALT_INV_RegFile[30][20]~q\,
	datad => \ALT_INV_RegFile[29][20]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux70~22_combout\,
	datag => \ALT_INV_RegFile[28][20]~q\,
	combout => \Mux70~9_combout\);

-- Location: FF_X60_Y1_N52
\RegFile[18][20]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][20]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][20]~DUPLICATE_q\);

-- Location: MLABCELL_X65_Y2_N0
\Mux70~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux70~18_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[16][20]~q\))) # (\R.curInst\(15) & (\RegFile[17][20]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[18][20]~DUPLICATE_q\))) # (\R.curInst\(15) & (\RegFile[19][20]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[19][20]~q\,
	datab => \ALT_INV_RegFile[17][20]~q\,
	datac => \ALT_INV_RegFile[18][20]~DUPLICATE_q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][20]~q\,
	combout => \Mux70~18_combout\);

-- Location: MLABCELL_X65_Y2_N48
\Mux70~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux70~5_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux70~18_combout\)))) # (\R.curInst\(17) & ((!\Mux70~18_combout\ & ((\RegFile[20][20]~q\))) # (\Mux70~18_combout\ & (\RegFile[21][20]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux70~18_combout\)))) # (\R.curInst\(17) & ((!\Mux70~18_combout\ & ((\RegFile[22][20]~q\))) # (\Mux70~18_combout\ & (\RegFile[23][20]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[23][20]~q\,
	datab => \ALT_INV_RegFile[21][20]~q\,
	datac => \ALT_INV_RegFile[22][20]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux70~18_combout\,
	datag => \ALT_INV_RegFile[20][20]~q\,
	combout => \Mux70~5_combout\);

-- Location: LABCELL_X67_Y3_N21
\Mux70~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux70~13_combout\ = ( \Mux70~9_combout\ & ( \Mux70~5_combout\ & ( ((!\R.curInst\(18) & (\Mux70~26_combout\)) # (\R.curInst\(18) & ((\Mux70~1_combout\)))) # (\R.curInst\(19)) ) ) ) # ( !\Mux70~9_combout\ & ( \Mux70~5_combout\ & ( (!\R.curInst\(18) & 
-- (((\R.curInst\(19))) # (\Mux70~26_combout\))) # (\R.curInst\(18) & (((\Mux70~1_combout\ & !\R.curInst\(19))))) ) ) ) # ( \Mux70~9_combout\ & ( !\Mux70~5_combout\ & ( (!\R.curInst\(18) & (\Mux70~26_combout\ & ((!\R.curInst\(19))))) # (\R.curInst\(18) & 
-- (((\R.curInst\(19)) # (\Mux70~1_combout\)))) ) ) ) # ( !\Mux70~9_combout\ & ( !\Mux70~5_combout\ & ( (!\R.curInst\(19) & ((!\R.curInst\(18) & (\Mux70~26_combout\)) # (\R.curInst\(18) & ((\Mux70~1_combout\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010011100000000001001110101010100100111101010100010011111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(18),
	datab => \ALT_INV_Mux70~26_combout\,
	datac => \ALT_INV_Mux70~1_combout\,
	datad => \ALT_INV_R.curInst\(19),
	datae => \ALT_INV_Mux70~9_combout\,
	dataf => \ALT_INV_Mux70~5_combout\,
	combout => \Mux70~13_combout\);

-- Location: LABCELL_X73_Y5_N3
\Mux234~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux234~0_combout\ = ( \Mux70~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC\(20)))) ) ) # ( !\Mux70~13_combout\ & ( (\vAluSrc1~2_combout\ & (!\vAluSrc1~1_combout\ & \R.curPC\(20))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010000000000000101000010100000111100001010000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluSrc1~2_combout\,
	datac => \ALT_INV_vAluSrc1~1_combout\,
	datad => \ALT_INV_R.curPC\(20),
	dataf => \ALT_INV_Mux70~13_combout\,
	combout => \Mux234~0_combout\);

-- Location: LABCELL_X74_Y5_N18
\ShiftLeft0~36\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~36_combout\ = ( \NxR.aluData2[1]~17_combout\ & ( \Mux232~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (\Mux234~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & ((\Mux235~0_combout\))) ) ) ) # ( !\NxR.aluData2[1]~17_combout\ & ( 
-- \Mux232~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\) # (\Mux233~0_combout\) ) ) ) # ( \NxR.aluData2[1]~17_combout\ & ( !\Mux232~0_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (\Mux234~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & 
-- ((\Mux235~0_combout\))) ) ) ) # ( !\NxR.aluData2[1]~17_combout\ & ( !\Mux232~0_combout\ & ( (\Mux233~0_combout\ & \NxR.aluData2[0]~16_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101001100000011111111110101111101010011000000111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux233~0_combout\,
	datab => \ALT_INV_Mux234~0_combout\,
	datac => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datad => \ALT_INV_Mux235~0_combout\,
	datae => \ALT_INV_NxR.aluData2[1]~17_combout\,
	dataf => \ALT_INV_Mux232~0_combout\,
	combout => \ShiftLeft0~36_combout\);

-- Location: FF_X74_Y5_N19
\ShiftLeft0~36_NEW_REG602\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~36_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~36_OTERM603\);

-- Location: LABCELL_X74_Y3_N24
\ShiftLeft0~45\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~45_combout\ = ( \NxR.aluData2[0]~16_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( \Mux231~0_combout\ ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( \Mux230~0_combout\ ) ) ) # ( \NxR.aluData2[0]~16_combout\ & ( 
-- !\NxR.aluData2[1]~17_combout\ & ( \Mux229~0_combout\ ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( !\NxR.aluData2[1]~17_combout\ & ( \Mux228~0_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111000011110000111101010101010101010011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux230~0_combout\,
	datab => \ALT_INV_Mux231~0_combout\,
	datac => \ALT_INV_Mux229~0_combout\,
	datad => \ALT_INV_Mux228~0_combout\,
	datae => \ALT_INV_NxR.aluData2[0]~16_combout\,
	dataf => \ALT_INV_NxR.aluData2[1]~17_combout\,
	combout => \ShiftLeft0~45_combout\);

-- Location: FF_X74_Y3_N25
\ShiftLeft0~45_NEW_REG756\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~45_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~45_OTERM757\);

-- Location: LABCELL_X73_Y5_N6
\ShiftLeft0~53\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~53_combout\ = ( \Mux227~0_combout\ & ( \NxR.aluData2[0]~16_combout\ & ( (\NxR.aluData2[1]~17_combout\) # (\Mux225~0_combout\) ) ) ) # ( !\Mux227~0_combout\ & ( \NxR.aluData2[0]~16_combout\ & ( (\Mux225~0_combout\ & 
-- !\NxR.aluData2[1]~17_combout\) ) ) ) # ( \Mux227~0_combout\ & ( !\NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (\Mux224~0_combout\)) # (\NxR.aluData2[1]~17_combout\ & ((\Mux226~0_combout\))) ) ) ) # ( !\Mux227~0_combout\ & ( 
-- !\NxR.aluData2[0]~16_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (\Mux224~0_combout\)) # (\NxR.aluData2[1]~17_combout\ & ((\Mux226~0_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100001111001100110000111101010101000000000101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux225~0_combout\,
	datab => \ALT_INV_Mux224~0_combout\,
	datac => \ALT_INV_Mux226~0_combout\,
	datad => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datae => \ALT_INV_Mux227~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[0]~16_combout\,
	combout => \ShiftLeft0~53_combout\);

-- Location: FF_X73_Y5_N7
\ShiftLeft0~53_NEW_REG764\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~53_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~53_OTERM765\);

-- Location: MLABCELL_X78_Y7_N30
\ShiftLeft0~54\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~54_combout\ = ( \ShiftLeft0~53_OTERM765\ & ( \R.aluData2\(3) & ( (!\R.aluData2\(2) & (\ShiftLeft0~36_OTERM603\)) # (\R.aluData2\(2) & ((\ShiftLeft0~28_OTERM295\))) ) ) ) # ( !\ShiftLeft0~53_OTERM765\ & ( \R.aluData2\(3) & ( (!\R.aluData2\(2) & 
-- (\ShiftLeft0~36_OTERM603\)) # (\R.aluData2\(2) & ((\ShiftLeft0~28_OTERM295\))) ) ) ) # ( \ShiftLeft0~53_OTERM765\ & ( !\R.aluData2\(3) & ( (!\R.aluData2\(2)) # (\ShiftLeft0~45_OTERM757\) ) ) ) # ( !\ShiftLeft0~53_OTERM765\ & ( !\R.aluData2\(3) & ( 
-- (\ShiftLeft0~45_OTERM757\ & \R.aluData2\(2)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110011111111110011001101010101000011110101010100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~36_OTERM603\,
	datab => \ALT_INV_ShiftLeft0~45_OTERM757\,
	datac => \ALT_INV_ShiftLeft0~28_OTERM295\,
	datad => \ALT_INV_R.aluData2\(2),
	datae => \ALT_INV_ShiftLeft0~53_OTERM765\,
	dataf => \ALT_INV_R.aluData2\(3),
	combout => \ShiftLeft0~54_combout\);

-- Location: MLABCELL_X72_Y6_N54
\Selector2~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector2~0_combout\ = ( \R.aluOp.ALUOpSRL~q\ & ( \R.aluOp.ALUOpSRA~q\ & ( (!\ShiftRight0~7_OTERM233DUPLICATE_q\ & (((\ShiftRight1~28_OTERM23\)) # (\ShiftRight0~2_OTERM25\))) # (\ShiftRight0~7_OTERM233DUPLICATE_q\ & (((\R.aluData1\(31))))) ) ) ) # ( 
-- !\R.aluOp.ALUOpSRL~q\ & ( \R.aluOp.ALUOpSRA~q\ & ( (!\ShiftRight0~7_OTERM233DUPLICATE_q\ & ((\ShiftRight1~28_OTERM23\))) # (\ShiftRight0~7_OTERM233DUPLICATE_q\ & (\R.aluData1\(31))) ) ) ) # ( \R.aluOp.ALUOpSRL~q\ & ( !\R.aluOp.ALUOpSRA~q\ & ( 
-- (!\ShiftRight0~7_OTERM233DUPLICATE_q\ & \ShiftRight0~2_OTERM25\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000001000100010001000000101101011110010011110101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight0~7_OTERM233DUPLICATE_q\,
	datab => \ALT_INV_ShiftRight0~2_OTERM25\,
	datac => \ALT_INV_R.aluData1\(31),
	datad => \ALT_INV_ShiftRight1~28_OTERM23\,
	datae => \ALT_INV_R.aluOp.ALUOpSRL~q\,
	dataf => \ALT_INV_R.aluOp.ALUOpSRA~q\,
	combout => \Selector2~0_combout\);

-- Location: LABCELL_X79_Y7_N0
\Selector2~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector2~1_combout\ = ( !\Selector17~0_OTERM391\ & ( \R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( (!\R.aluData1\(30) & ((!\R.aluData2\(30)) # ((!\R.aluOp.ALUOpOr~q\ & !\R.aluOp.ALUOpXor~DUPLICATE_q\)))) # (\R.aluData1\(30) & (!\R.aluOp.ALUOpOr~q\ & 
-- (!\R.aluOp.ALUOpXor~DUPLICATE_q\ & !\R.aluData2\(30)))) ) ) ) # ( !\Selector17~0_OTERM391\ & ( !\R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( (!\R.aluOp.ALUOpOr~q\ & ((!\R.aluOp.ALUOpXor~DUPLICATE_q\) # (!\R.aluData1\(30) $ (\R.aluData2\(30))))) # 
-- (\R.aluOp.ALUOpOr~q\ & (((!\R.aluData1\(30) & !\R.aluData2\(30))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111100010001010000000000000000011111000100000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpOr~q\,
	datab => \ALT_INV_R.aluOp.ALUOpXor~DUPLICATE_q\,
	datac => \ALT_INV_R.aluData1\(30),
	datad => \ALT_INV_R.aluData2\(30),
	datae => \ALT_INV_Selector17~0_OTERM391\,
	dataf => \ALT_INV_R.aluOp.ALUOpAnd~DUPLICATE_q\,
	combout => \Selector2~1_combout\);

-- Location: LABCELL_X77_Y7_N6
\Selector2~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector2~2_combout\ = ( \Selector2~1_combout\ & ( \R.aluData2\(4) & ( (\ShiftLeft0~21_combout\ & \R.aluOp.ALUOpSLL~q\) ) ) ) # ( !\Selector2~1_combout\ & ( \R.aluData2\(4) ) ) # ( \Selector2~1_combout\ & ( !\R.aluData2\(4) & ( ((\ShiftLeft0~54_combout\ 
-- & \R.aluOp.ALUOpSLL~q\)) # (\Selector2~0_combout\) ) ) ) # ( !\Selector2~1_combout\ & ( !\R.aluData2\(4) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111001100110111011111111111111111110000000000001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~54_combout\,
	datab => \ALT_INV_Selector2~0_combout\,
	datac => \ALT_INV_ShiftLeft0~21_combout\,
	datad => \ALT_INV_R.aluOp.ALUOpSLL~q\,
	datae => \ALT_INV_Selector2~1_combout\,
	dataf => \ALT_INV_R.aluData2\(4),
	combout => \Selector2~2_combout\);

-- Location: LABCELL_X77_Y3_N30
\Comb:vJumpAdr[30]~0_RESYN1036\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[30]~0_RESYN1036_BDD1037\ = ( \Add1~121_sumout\ & ( \Add2~121_sumout\ & ( (\R.aluOp.ALUOpAdd~q\) # (\R.aluOp.ALUOpSub~q\) ) ) ) # ( !\Add1~121_sumout\ & ( \Add2~121_sumout\ & ( \R.aluOp.ALUOpSub~q\ ) ) ) # ( \Add1~121_sumout\ & ( 
-- !\Add2~121_sumout\ & ( \R.aluOp.ALUOpAdd~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000111100110011001100110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datae => \ALT_INV_Add1~121_sumout\,
	dataf => \ALT_INV_Add2~121_sumout\,
	combout => \Comb:vJumpAdr[30]~0_RESYN1036_BDD1037\);

-- Location: FF_X77_Y3_N38
\R.curPC[30]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[30]~0_combout\,
	asdata => \Add0~113_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(30));

-- Location: LABCELL_X77_Y3_N0
\Add3~121\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~121_sumout\ = SUM(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux124~1_combout\)) ) + ( \R.curPC\(30) ) + ( \Add3~118\ ))
-- \Add3~122\ = CARRY(( (\R.curInst\(0) & (\R.curInst\(1) & \Mux124~1_combout\)) ) + ( \R.curPC\(30) ) + ( \Add3~118\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000010001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datac => \ALT_INV_R.curPC\(30),
	datad => \ALT_INV_Mux124~1_combout\,
	cin => \Add3~118\,
	sumout => \Add3~121_sumout\,
	cout => \Add3~122\);

-- Location: LABCELL_X77_Y3_N36
\Comb:vJumpAdr[30]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[30]~0_combout\ = ( \Add3~121_sumout\ & ( \R.aluRes\(30) & ( (((!\Equal4~2_combout\) # (!\R.aluCalc~q\)) # (\Comb:vJumpAdr[30]~0_RESYN1036_BDD1037\)) # (\Selector2~2_combout\) ) ) ) # ( !\Add3~121_sumout\ & ( \R.aluRes\(30) & ( 
-- (\Equal4~2_combout\ & (((!\R.aluCalc~q\) # (\Comb:vJumpAdr[30]~0_RESYN1036_BDD1037\)) # (\Selector2~2_combout\))) ) ) ) # ( \Add3~121_sumout\ & ( !\R.aluRes\(30) & ( (!\Equal4~2_combout\) # ((\R.aluCalc~q\ & ((\Comb:vJumpAdr[30]~0_RESYN1036_BDD1037\) # 
-- (\Selector2~2_combout\)))) ) ) ) # ( !\Add3~121_sumout\ & ( !\R.aluRes\(30) & ( (\Equal4~2_combout\ & (\R.aluCalc~q\ & ((\Comb:vJumpAdr[30]~0_RESYN1036_BDD1037\) # (\Selector2~2_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000111111100001111011100001111000001111111111111110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector2~2_combout\,
	datab => \ALT_INV_Comb:vJumpAdr[30]~0_RESYN1036_BDD1037\,
	datac => \ALT_INV_Equal4~2_combout\,
	datad => \ALT_INV_R.aluCalc~q\,
	datae => \ALT_INV_Add3~121_sumout\,
	dataf => \ALT_INV_R.aluRes\(30),
	combout => \Comb:vJumpAdr[30]~0_combout\);

-- Location: FF_X77_Y3_N37
\R.curPC[30]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[30]~0_combout\,
	asdata => \Add0~113_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC[30]~DUPLICATE_q\);

-- Location: LABCELL_X81_Y5_N57
\Add0~117\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~117_sumout\ = SUM(( GND ) + ( GND ) + ( \Add0~114\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	cin => \Add0~114\,
	sumout => \Add0~117_sumout\);

-- Location: IOIBUF_X22_Y0_N1
\avm_d_readdata[7]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(7),
	o => \avm_d_readdata[7]~input_o\);

-- Location: LABCELL_X79_Y2_N33
\Comb:vRegWriteData[31]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[31]~1_combout\ = ( \avm_d_readdata[23]~input_o\ & ( \avm_d_readdata[7]~input_o\ & ( (!\R.curInst\(14) & ((!\R.curInst\(12) & ((\R.curInst\(13)) # (\avm_d_readdata[31]~input_o\))) # (\R.curInst\(12) & ((!\R.curInst\(13)))))) ) ) ) # ( 
-- !\avm_d_readdata[23]~input_o\ & ( \avm_d_readdata[7]~input_o\ & ( (!\R.curInst\(12) & (!\R.curInst\(14) & ((\R.curInst\(13)) # (\avm_d_readdata[31]~input_o\)))) ) ) ) # ( \avm_d_readdata[23]~input_o\ & ( !\avm_d_readdata[7]~input_o\ & ( (!\R.curInst\(14) 
-- & (!\R.curInst\(13) & ((\avm_d_readdata[31]~input_o\) # (\R.curInst\(12))))) ) ) ) # ( !\avm_d_readdata[23]~input_o\ & ( !\avm_d_readdata[7]~input_o\ & ( (!\R.curInst\(12) & (\avm_d_readdata[31]~input_o\ & (!\R.curInst\(14) & !\R.curInst\(13)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010000000000000011100000000000000100000101000000111000010100000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(12),
	datab => \ALT_INV_avm_d_readdata[31]~input_o\,
	datac => \ALT_INV_R.curInst\(14),
	datad => \ALT_INV_R.curInst\(13),
	datae => \ALT_INV_avm_d_readdata[23]~input_o\,
	dataf => \ALT_INV_avm_d_readdata[7]~input_o\,
	combout => \Comb:vRegWriteData[31]~1_combout\);

-- Location: MLABCELL_X78_Y5_N48
\Comb:vRegWriteData[31]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[31]~2_combout\ = ( \Comb:vRegWriteData[31]~1_combout\ & ( (!\R.memToReg~q\ & (!\Selector1~2_combout\ & ((!\R.aluOp.ALUOpAdd~q\) # (!\Add1~125_sumout\)))) ) ) # ( !\Comb:vRegWriteData[31]~1_combout\ & ( ((!\Selector1~2_combout\ & 
-- ((!\R.aluOp.ALUOpAdd~q\) # (!\Add1~125_sumout\)))) # (\R.memToReg~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111110101010101111111010101010110101000000000001010100000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.memToReg~q\,
	datab => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datac => \ALT_INV_Add1~125_sumout\,
	datad => \ALT_INV_Selector1~2_combout\,
	dataf => \ALT_INV_Comb:vRegWriteData[31]~1_combout\,
	combout => \Comb:vRegWriteData[31]~2_combout\);

-- Location: MLABCELL_X78_Y5_N42
\Comb:vRegWriteData[31]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[31]~0_combout\ = ( \Add2~125_sumout\ & ( \Comb:vRegWriteData[31]~2_combout\ & ( (!\R.memToReg~q\ & ((!\R.aluCalc~q\ & ((\R.aluRes\(31)))) # (\R.aluCalc~q\ & (\R.aluOp.ALUOpSub~q\)))) ) ) ) # ( !\Add2~125_sumout\ & ( 
-- \Comb:vRegWriteData[31]~2_combout\ & ( (!\R.aluCalc~q\ & (!\R.memToReg~q\ & \R.aluRes\(31))) ) ) ) # ( \Add2~125_sumout\ & ( !\Comb:vRegWriteData[31]~2_combout\ & ( ((\R.aluRes\(31)) # (\R.memToReg~q\)) # (\R.aluCalc~q\) ) ) ) # ( !\Add2~125_sumout\ & ( 
-- !\Comb:vRegWriteData[31]~2_combout\ & ( ((\R.aluRes\(31)) # (\R.memToReg~q\)) # (\R.aluCalc~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101111111111111010111111111111100000000101000000001000010110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluCalc~q\,
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_R.memToReg~q\,
	datad => \ALT_INV_R.aluRes\(31),
	datae => \ALT_INV_Add2~125_sumout\,
	dataf => \ALT_INV_Comb:vRegWriteData[31]~2_combout\,
	combout => \Comb:vRegWriteData[31]~0_combout\);

-- Location: FF_X81_Y5_N59
\R.regWriteData[31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Add0~117_sumout\,
	asdata => \Comb:vRegWriteData[31]~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(31));

-- Location: FF_X68_Y5_N14
\RegFile[3][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(31),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][31]~q\);

-- Location: FF_X70_Y5_N13
\RegFile[2][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(31),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][31]~q\);

-- Location: FF_X70_Y5_N19
\RegFile[7][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(31),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][31]~q\);

-- Location: FF_X59_Y4_N13
\RegFile[5][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(31),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][31]~q\);

-- Location: LABCELL_X67_Y5_N24
\RegFile[4][31]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[4][31]~feeder_combout\ = ( \R.regWriteData\(31) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(31),
	combout => \RegFile[4][31]~feeder_combout\);

-- Location: FF_X67_Y5_N25
\RegFile[4][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[4][31]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][31]~q\);

-- Location: FF_X68_Y5_N43
\RegFile[6][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(31),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][31]~q\);

-- Location: LABCELL_X68_Y5_N42
\Mux91~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux91~0_combout\ = ( \RegFile[6][31]~q\ & ( \R.curInst\(20) & ( (!\R.curInst\(21) & ((\RegFile[5][31]~q\))) # (\R.curInst\(21) & (\RegFile[7][31]~q\)) ) ) ) # ( !\RegFile[6][31]~q\ & ( \R.curInst\(20) & ( (!\R.curInst\(21) & ((\RegFile[5][31]~q\))) # 
-- (\R.curInst\(21) & (\RegFile[7][31]~q\)) ) ) ) # ( \RegFile[6][31]~q\ & ( !\R.curInst\(20) & ( (\R.curInst\(21)) # (\RegFile[4][31]~q\) ) ) ) # ( !\RegFile[6][31]~q\ & ( !\R.curInst\(20) & ( (\RegFile[4][31]~q\ & !\R.curInst\(21)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100000000000011111111111100110011010101010011001101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[7][31]~q\,
	datab => \ALT_INV_RegFile[5][31]~q\,
	datac => \ALT_INV_RegFile[4][31]~q\,
	datad => \ALT_INV_R.curInst\(21),
	datae => \ALT_INV_RegFile[6][31]~q\,
	dataf => \ALT_INV_R.curInst\(20),
	combout => \Mux91~0_combout\);

-- Location: MLABCELL_X72_Y3_N36
\RegFile[1][31]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[1][31]~feeder_combout\ = \R.regWriteData\(31)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.regWriteData\(31),
	combout => \RegFile[1][31]~feeder_combout\);

-- Location: FF_X72_Y3_N37
\RegFile[1][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[1][31]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][31]~q\);

-- Location: LABCELL_X68_Y5_N12
\Mux91~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux91~26_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (\RegFile[1][31]~q\ & (\R.curInst\(20)))) # (\R.curInst\(22) & (((\Mux91~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (((\RegFile[2][31]~q\)))) # 
-- (\R.curInst\(20) & (\RegFile[3][31]~q\)))) # (\R.curInst\(22) & ((((\Mux91~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001100000011000100010000110011001111110011111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][31]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[2][31]~q\,
	datad => \ALT_INV_R.curInst\(20),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux91~0_combout\,
	datag => \ALT_INV_RegFile[1][31]~q\,
	combout => \Mux91~26_combout\);

-- Location: FF_X65_Y1_N44
\RegFile[13][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(31),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][31]~q\);

-- Location: FF_X66_Y1_N32
\RegFile[15][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(31),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][31]~q\);

-- Location: LABCELL_X66_Y1_N0
\RegFile[14][31]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[14][31]~feeder_combout\ = ( \R.regWriteData\(31) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(31),
	combout => \RegFile[14][31]~feeder_combout\);

-- Location: FF_X66_Y1_N2
\RegFile[14][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[14][31]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][31]~q\);

-- Location: FF_X66_Y1_N44
\RegFile[9][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(31),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][31]~q\);

-- Location: FF_X65_Y1_N8
\RegFile[11][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(31),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][31]~q\);

-- Location: LABCELL_X61_Y1_N18
\RegFile[10][31]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[10][31]~feeder_combout\ = ( \R.regWriteData\(31) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(31),
	combout => \RegFile[10][31]~feeder_combout\);

-- Location: FF_X61_Y1_N19
\RegFile[10][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[10][31]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][31]~q\);

-- Location: FF_X59_Y1_N1
\RegFile[8][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(31),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][31]~q\);

-- Location: LABCELL_X66_Y1_N42
\Mux91~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux91~14_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[8][31]~q\))) # (\R.curInst\(20) & (\RegFile[9][31]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[10][31]~q\))) # (\R.curInst\(20) & (\RegFile[11][31]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][31]~q\,
	datab => \ALT_INV_RegFile[11][31]~q\,
	datac => \ALT_INV_RegFile[10][31]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][31]~q\,
	combout => \Mux91~14_combout\);

-- Location: LABCELL_X74_Y1_N36
\RegFile[12][31]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[12][31]~feeder_combout\ = ( \R.regWriteData\(31) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(31),
	combout => \RegFile[12][31]~feeder_combout\);

-- Location: FF_X74_Y1_N37
\RegFile[12][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[12][31]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][31]~q\);

-- Location: LABCELL_X66_Y1_N30
\Mux91~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux91~1_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux91~14_combout\)))) # (\R.curInst\(22) & ((!\Mux91~14_combout\ & ((\RegFile[12][31]~q\))) # (\Mux91~14_combout\ & (\RegFile[13][31]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux91~14_combout\)))) # (\R.curInst\(22) & ((!\Mux91~14_combout\ & ((\RegFile[14][31]~q\))) # (\Mux91~14_combout\ & (\RegFile[15][31]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][31]~q\,
	datab => \ALT_INV_RegFile[15][31]~q\,
	datac => \ALT_INV_RegFile[14][31]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux91~14_combout\,
	datag => \ALT_INV_RegFile[12][31]~q\,
	combout => \Mux91~1_combout\);

-- Location: FF_X72_Y6_N50
\RegFile[29][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(31),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][31]~q\);

-- Location: FF_X57_Y6_N52
\RegFile[30][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(31),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][31]~q\);

-- Location: FF_X65_Y4_N26
\RegFile[31][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(31),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][31]~q\);

-- Location: FF_X65_Y4_N56
\RegFile[25][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(31),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][31]~q\);

-- Location: FF_X65_Y4_N14
\RegFile[27][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(31),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][31]~q\);

-- Location: FF_X67_Y4_N1
\RegFile[26][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(31),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][31]~q\);

-- Location: LABCELL_X57_Y4_N45
\RegFile[24][31]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[24][31]~feeder_combout\ = ( \R.regWriteData\(31) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(31),
	combout => \RegFile[24][31]~feeder_combout\);

-- Location: FF_X57_Y4_N46
\RegFile[24][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[24][31]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][31]~q\);

-- Location: MLABCELL_X65_Y4_N54
\Mux91~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux91~22_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[24][31]~q\))) # (\R.curInst\(20) & (\RegFile[25][31]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[26][31]~q\))) # (\R.curInst\(20) & (\RegFile[27][31]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[25][31]~q\,
	datab => \ALT_INV_RegFile[27][31]~q\,
	datac => \ALT_INV_RegFile[26][31]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][31]~q\,
	combout => \Mux91~22_combout\);

-- Location: LABCELL_X71_Y8_N9
\RegFile[28][31]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[28][31]~feeder_combout\ = ( \R.regWriteData\(31) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(31),
	combout => \RegFile[28][31]~feeder_combout\);

-- Location: FF_X71_Y8_N11
\RegFile[28][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[28][31]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][31]~q\);

-- Location: MLABCELL_X72_Y6_N48
\Mux91~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux91~9_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux91~22_combout\))))) # (\R.curInst\(22) & (((!\Mux91~22_combout\ & ((\RegFile[28][31]~q\))) # (\Mux91~22_combout\ & (\RegFile[29][31]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux91~22_combout\)))) # (\R.curInst\(22) & ((!\Mux91~22_combout\ & (\RegFile[30][31]~q\)) # (\Mux91~22_combout\ & ((\RegFile[31][31]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[29][31]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[30][31]~q\,
	datad => \ALT_INV_RegFile[31][31]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux91~22_combout\,
	datag => \ALT_INV_RegFile[28][31]~q\,
	combout => \Mux91~9_combout\);

-- Location: FF_X72_Y4_N50
\RegFile[21][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(31),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][31]~q\);

-- Location: FF_X70_Y5_N49
\RegFile[23][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(31),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][31]~q\);

-- Location: LABCELL_X61_Y8_N51
\RegFile[22][31]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[22][31]~feeder_combout\ = ( \R.regWriteData\(31) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(31),
	combout => \RegFile[22][31]~feeder_combout\);

-- Location: FF_X61_Y8_N52
\RegFile[22][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[22][31]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][31]~q\);

-- Location: FF_X66_Y4_N2
\RegFile[17][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(31),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][31]~q\);

-- Location: LABCELL_X66_Y4_N24
\RegFile[18][31]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[18][31]~feeder_combout\ = ( \R.regWriteData\(31) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(31),
	combout => \RegFile[18][31]~feeder_combout\);

-- Location: FF_X66_Y4_N26
\RegFile[18][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][31]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][31]~q\);

-- Location: LABCELL_X66_Y4_N54
\RegFile[19][31]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[19][31]~feeder_combout\ = ( \R.regWriteData\(31) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(31),
	combout => \RegFile[19][31]~feeder_combout\);

-- Location: FF_X66_Y4_N55
\RegFile[19][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[19][31]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][31]~q\);

-- Location: LABCELL_X61_Y8_N24
\RegFile[16][31]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[16][31]~feeder_combout\ = ( \R.regWriteData\(31) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(31),
	combout => \RegFile[16][31]~feeder_combout\);

-- Location: FF_X61_Y8_N25
\RegFile[16][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[16][31]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][31]~q\);

-- Location: LABCELL_X66_Y4_N0
\Mux91~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux91~18_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[16][31]~q\))) # (\R.curInst\(20) & (\RegFile[17][31]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & (\RegFile[18][31]~q\)) # (\R.curInst\(20) & ((\RegFile[19][31]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[17][31]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[18][31]~q\,
	datad => \ALT_INV_RegFile[19][31]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][31]~q\,
	combout => \Mux91~18_combout\);

-- Location: LABCELL_X68_Y6_N21
\RegFile[20][31]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[20][31]~feeder_combout\ = ( \R.regWriteData\(31) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(31),
	combout => \RegFile[20][31]~feeder_combout\);

-- Location: FF_X68_Y6_N22
\RegFile[20][31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[20][31]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][31]~q\);

-- Location: MLABCELL_X72_Y4_N48
\Mux91~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux91~5_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux91~18_combout\)))) # (\R.curInst\(22) & ((!\Mux91~18_combout\ & ((\RegFile[20][31]~q\))) # (\Mux91~18_combout\ & (\RegFile[21][31]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux91~18_combout\)))) # (\R.curInst\(22) & ((!\Mux91~18_combout\ & ((\RegFile[22][31]~q\))) # (\Mux91~18_combout\ & (\RegFile[23][31]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][31]~q\,
	datab => \ALT_INV_RegFile[23][31]~q\,
	datac => \ALT_INV_RegFile[22][31]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux91~18_combout\,
	datag => \ALT_INV_RegFile[20][31]~q\,
	combout => \Mux91~5_combout\);

-- Location: MLABCELL_X72_Y5_N30
\Mux91~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux91~13_combout\ = ( \Mux91~9_combout\ & ( \Mux91~5_combout\ & ( ((!\R.curInst\(23) & (\Mux91~26_combout\)) # (\R.curInst\(23) & ((\Mux91~1_combout\)))) # (\R.curInst\(24)) ) ) ) # ( !\Mux91~9_combout\ & ( \Mux91~5_combout\ & ( (!\R.curInst\(23) & 
-- (((\Mux91~26_combout\)) # (\R.curInst\(24)))) # (\R.curInst\(23) & (!\R.curInst\(24) & ((\Mux91~1_combout\)))) ) ) ) # ( \Mux91~9_combout\ & ( !\Mux91~5_combout\ & ( (!\R.curInst\(23) & (!\R.curInst\(24) & (\Mux91~26_combout\))) # (\R.curInst\(23) & 
-- (((\Mux91~1_combout\)) # (\R.curInst\(24)))) ) ) ) # ( !\Mux91~9_combout\ & ( !\Mux91~5_combout\ & ( (!\R.curInst\(24) & ((!\R.curInst\(23) & (\Mux91~26_combout\)) # (\R.curInst\(23) & ((\Mux91~1_combout\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000100001001100000110010101110100101010011011100011101101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(23),
	datab => \ALT_INV_R.curInst\(24),
	datac => \ALT_INV_Mux91~26_combout\,
	datad => \ALT_INV_Mux91~1_combout\,
	datae => \ALT_INV_Mux91~9_combout\,
	dataf => \ALT_INV_Mux91~5_combout\,
	combout => \Mux91~13_combout\);

-- Location: MLABCELL_X72_Y5_N45
\NxR.aluData2[31]~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[31]~29_combout\ = ( \Mux91~13_combout\ & ( (!\vAluSrc2~1_combout\) # ((\Mux123~3_combout\ & \Equal4~1_combout\)) ) ) # ( !\Mux91~13_combout\ & ( (\Mux123~3_combout\ & (\Equal4~1_combout\ & \vAluSrc2~1_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000011000000000000001111111111000000111111111100000011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Mux123~3_combout\,
	datac => \ALT_INV_Equal4~1_combout\,
	datad => \ALT_INV_vAluSrc2~1_combout\,
	dataf => \ALT_INV_Mux91~13_combout\,
	combout => \NxR.aluData2[31]~29_combout\);

-- Location: FF_X72_Y5_N23
\R.aluData2[31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \NxR.aluData2[31]~29_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData2\(31));

-- Location: MLABCELL_X82_Y5_N36
\Selector1~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector1~3_combout\ = ( \Add1~125_sumout\ & ( (((\Add2~125_sumout\ & \R.aluOp.ALUOpSub~q\)) # (\Selector1~2_combout\)) # (\R.aluOp.ALUOpAdd~q\) ) ) # ( !\Add1~125_sumout\ & ( ((\Add2~125_sumout\ & \R.aluOp.ALUOpSub~q\)) # (\Selector1~2_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000111111111000100011111111100011111111111110001111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add2~125_sumout\,
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_Selector1~2_combout\,
	dataf => \ALT_INV_Add1~125_sumout\,
	combout => \Selector1~3_combout\);

-- Location: FF_X82_Y5_N37
\R.aluRes[31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector1~3_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(31));

-- Location: LABCELL_X77_Y3_N6
\vAluRes~30\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~30_combout\ = ( !\R.aluCalc~q\ & ( \R.aluRes\(31) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluRes\(31),
	dataf => \ALT_INV_R.aluCalc~q\,
	combout => \vAluRes~30_combout\);

-- Location: LABCELL_X77_Y3_N24
\vAluRes~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~29_combout\ = ( \Add1~125_sumout\ & ( \Selector1~2_combout\ & ( \R.aluCalc~q\ ) ) ) # ( !\Add1~125_sumout\ & ( \Selector1~2_combout\ & ( \R.aluCalc~q\ ) ) ) # ( \Add1~125_sumout\ & ( !\Selector1~2_combout\ & ( (\R.aluCalc~q\ & 
-- (((\R.aluOp.ALUOpSub~q\ & \Add2~125_sumout\)) # (\R.aluOp.ALUOpAdd~q\))) ) ) ) # ( !\Add1~125_sumout\ & ( !\Selector1~2_combout\ & ( (\R.aluCalc~q\ & (\R.aluOp.ALUOpSub~q\ & \Add2~125_sumout\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000010001000001010001010101010101010101010101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluCalc~q\,
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_Add2~125_sumout\,
	datae => \ALT_INV_Add1~125_sumout\,
	dataf => \ALT_INV_Selector1~2_combout\,
	combout => \vAluRes~29_combout\);

-- Location: FF_X77_Y3_N56
\R.curPC[31]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[31]~0_combout\,
	asdata => \Add0~117_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(31));

-- Location: LABCELL_X77_Y3_N3
\Add3~125\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add3~125_sumout\ = SUM(( \R.curPC\(31) ) + ( (\R.curInst\(0) & (\R.curInst\(1) & \Mux123~3_combout\)) ) + ( \Add3~122\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111101111111000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(0),
	datab => \ALT_INV_R.curInst\(1),
	datac => \ALT_INV_Mux123~3_combout\,
	datad => \ALT_INV_R.curPC\(31),
	cin => \Add3~122\,
	sumout => \Add3~125_sumout\);

-- Location: LABCELL_X77_Y3_N54
\Comb:vJumpAdr[31]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[31]~0_combout\ = ( \Add3~125_sumout\ & ( (!\Equal4~2_combout\) # ((\vAluRes~29_combout\) # (\vAluRes~30_combout\)) ) ) # ( !\Add3~125_sumout\ & ( (\Equal4~2_combout\ & ((\vAluRes~29_combout\) # (\vAluRes~30_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001010100010101101111111011111100010101000101011011111110111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Equal4~2_combout\,
	datab => \ALT_INV_vAluRes~30_combout\,
	datac => \ALT_INV_vAluRes~29_combout\,
	datae => \ALT_INV_Add3~125_sumout\,
	combout => \Comb:vJumpAdr[31]~0_combout\);

-- Location: FF_X77_Y3_N55
\R.curPC[31]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[31]~0_combout\,
	asdata => \Add0~117_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC[31]~DUPLICATE_q\);

-- Location: LABCELL_X71_Y5_N33
\Mux59~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux59~0_combout\ = ( \R.curInst\(15) & ( \R.curInst\(16) & ( \RegFile[7][31]~q\ ) ) ) # ( !\R.curInst\(15) & ( \R.curInst\(16) & ( \RegFile[6][31]~q\ ) ) ) # ( \R.curInst\(15) & ( !\R.curInst\(16) & ( \RegFile[5][31]~q\ ) ) ) # ( !\R.curInst\(15) & ( 
-- !\R.curInst\(16) & ( \RegFile[4][31]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101001100110011001100000000111111110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[4][31]~q\,
	datab => \ALT_INV_RegFile[5][31]~q\,
	datac => \ALT_INV_RegFile[7][31]~q\,
	datad => \ALT_INV_RegFile[6][31]~q\,
	datae => \ALT_INV_R.curInst\(15),
	dataf => \ALT_INV_R.curInst\(16),
	combout => \Mux59~0_combout\);

-- Location: LABCELL_X71_Y5_N0
\Mux59~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux59~26_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (\R.curInst\(15) & (\RegFile[1][31]~q\))) # (\R.curInst\(17) & (((\Mux59~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & ((!\R.curInst\(15) & (((\RegFile[2][31]~q\)))) # 
-- (\R.curInst\(15) & (\RegFile[3][31]~q\)))) # (\R.curInst\(17) & ((((\Mux59~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000000000110110000000000000101111111110001101111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(15),
	datab => \ALT_INV_RegFile[3][31]~q\,
	datac => \ALT_INV_RegFile[2][31]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux59~0_combout\,
	datag => \ALT_INV_RegFile[1][31]~q\,
	combout => \Mux59~26_combout\);

-- Location: FF_X66_Y4_N25
\RegFile[18][31]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][31]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][31]~DUPLICATE_q\);

-- Location: LABCELL_X70_Y5_N54
\Mux59~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux59~18_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[16][31]~q\))) # (\R.curInst\(15) & (\RegFile[17][31]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[18][31]~DUPLICATE_q\))) # (\R.curInst\(15) & (\RegFile[19][31]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[17][31]~q\,
	datab => \ALT_INV_RegFile[19][31]~q\,
	datac => \ALT_INV_RegFile[18][31]~DUPLICATE_q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][31]~q\,
	combout => \Mux59~18_combout\);

-- Location: LABCELL_X71_Y5_N6
\Mux59~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux59~5_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux59~18_combout\)))) # (\R.curInst\(17) & ((!\Mux59~18_combout\ & ((\RegFile[20][31]~q\))) # (\Mux59~18_combout\ & (\RegFile[21][31]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux59~18_combout\)))) # (\R.curInst\(17) & ((!\Mux59~18_combout\ & ((\RegFile[22][31]~q\))) # (\Mux59~18_combout\ & (\RegFile[23][31]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][31]~q\,
	datab => \ALT_INV_RegFile[23][31]~q\,
	datac => \ALT_INV_RegFile[22][31]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux59~18_combout\,
	datag => \ALT_INV_RegFile[20][31]~q\,
	combout => \Mux59~5_combout\);

-- Location: MLABCELL_X65_Y1_N6
\Mux59~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux59~14_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[8][31]~q\))) # (\R.curInst\(15) & (\RegFile[9][31]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & (\RegFile[10][31]~q\)) # (\R.curInst\(15) & ((\RegFile[11][31]~q\))))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][31]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[10][31]~q\,
	datad => \ALT_INV_RegFile[11][31]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][31]~q\,
	combout => \Mux59~14_combout\);

-- Location: MLABCELL_X65_Y1_N42
\Mux59~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux59~1_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux59~14_combout\)))) # (\R.curInst\(17) & ((!\Mux59~14_combout\ & (\RegFile[12][31]~q\)) # (\Mux59~14_combout\ & ((\RegFile[13][31]~q\)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) 
-- & ((((\Mux59~14_combout\))))) # (\R.curInst\(17) & (((!\Mux59~14_combout\ & ((\RegFile[14][31]~q\))) # (\Mux59~14_combout\ & (\RegFile[15][31]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111001100111111111101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][31]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[14][31]~q\,
	datad => \ALT_INV_RegFile[13][31]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux59~14_combout\,
	datag => \ALT_INV_RegFile[12][31]~q\,
	combout => \Mux59~1_combout\);

-- Location: MLABCELL_X65_Y4_N12
\Mux59~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux59~22_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[24][31]~q\))) # (\R.curInst\(15) & (\RegFile[25][31]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[26][31]~q\))) # (\R.curInst\(15) & (\RegFile[27][31]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[25][31]~q\,
	datab => \ALT_INV_RegFile[27][31]~q\,
	datac => \ALT_INV_RegFile[26][31]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][31]~q\,
	combout => \Mux59~22_combout\);

-- Location: MLABCELL_X65_Y4_N24
\Mux59~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux59~9_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux59~22_combout\)))) # (\R.curInst\(17) & ((!\Mux59~22_combout\ & (\RegFile[28][31]~q\)) # (\Mux59~22_combout\ & ((\RegFile[29][31]~q\)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) 
-- & ((((\Mux59~22_combout\))))) # (\R.curInst\(17) & (((!\Mux59~22_combout\ & ((\RegFile[30][31]~q\))) # (\Mux59~22_combout\ & (\RegFile[31][31]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111001100111111111101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][31]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[30][31]~q\,
	datad => \ALT_INV_RegFile[29][31]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux59~22_combout\,
	datag => \ALT_INV_RegFile[28][31]~q\,
	combout => \Mux59~9_combout\);

-- Location: LABCELL_X71_Y5_N39
\Mux59~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux59~13_combout\ = ( \Mux59~1_combout\ & ( \Mux59~9_combout\ & ( ((!\R.curInst\(19) & (\Mux59~26_combout\)) # (\R.curInst\(19) & ((\Mux59~5_combout\)))) # (\R.curInst\(18)) ) ) ) # ( !\Mux59~1_combout\ & ( \Mux59~9_combout\ & ( (!\R.curInst\(18) & 
-- ((!\R.curInst\(19) & (\Mux59~26_combout\)) # (\R.curInst\(19) & ((\Mux59~5_combout\))))) # (\R.curInst\(18) & (((\R.curInst\(19))))) ) ) ) # ( \Mux59~1_combout\ & ( !\Mux59~9_combout\ & ( (!\R.curInst\(18) & ((!\R.curInst\(19) & (\Mux59~26_combout\)) # 
-- (\R.curInst\(19) & ((\Mux59~5_combout\))))) # (\R.curInst\(18) & (((!\R.curInst\(19))))) ) ) ) # ( !\Mux59~1_combout\ & ( !\Mux59~9_combout\ & ( (!\R.curInst\(18) & ((!\R.curInst\(19) & (\Mux59~26_combout\)) # (\R.curInst\(19) & ((\Mux59~5_combout\))))) ) 
-- ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100010000001100011101110000110001000100001111110111011100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux59~26_combout\,
	datab => \ALT_INV_R.curInst\(18),
	datac => \ALT_INV_Mux59~5_combout\,
	datad => \ALT_INV_R.curInst\(19),
	datae => \ALT_INV_Mux59~1_combout\,
	dataf => \ALT_INV_Mux59~9_combout\,
	combout => \Mux59~13_combout\);

-- Location: MLABCELL_X72_Y5_N57
\Mux223~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux223~0_combout\ = ( \Mux59~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC[31]~DUPLICATE_q\))) ) ) # ( !\Mux59~13_combout\ & ( (\R.curPC[31]~DUPLICATE_q\ & (\vAluSrc1~2_combout\ & !\vAluSrc1~1_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000000000000110000000011110011000000001111001100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.curPC[31]~DUPLICATE_q\,
	datac => \ALT_INV_vAluSrc1~2_combout\,
	datad => \ALT_INV_vAluSrc1~1_combout\,
	dataf => \ALT_INV_Mux59~13_combout\,
	combout => \Mux223~0_combout\);

-- Location: LABCELL_X71_Y7_N42
\ShiftRight1~48\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~48_combout\ = ( \Mux224~0_combout\ & ( \NxR.aluData2[2]~19_combout\ & ( ((!\NxR.aluData2[0]~16_combout\ & (!\NxR.aluData2[3]~18_combout\ & !\NxR.aluData2[1]~17_combout\))) # (\Mux223~0_combout\) ) ) ) # ( !\Mux224~0_combout\ & ( 
-- \NxR.aluData2[2]~19_combout\ & ( (\Mux223~0_combout\ & (((\NxR.aluData2[1]~17_combout\) # (\NxR.aluData2[3]~18_combout\)) # (\NxR.aluData2[0]~16_combout\))) ) ) ) # ( \Mux224~0_combout\ & ( !\NxR.aluData2[2]~19_combout\ & ( (\Mux223~0_combout\ & 
-- \NxR.aluData2[3]~18_combout\) ) ) ) # ( !\Mux224~0_combout\ & ( !\NxR.aluData2[2]~19_combout\ & ( (\Mux223~0_combout\ & \NxR.aluData2[3]~18_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101000001010000010100010101010101011101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux223~0_combout\,
	datab => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datac => \ALT_INV_NxR.aluData2[3]~18_combout\,
	datad => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datae => \ALT_INV_Mux224~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[2]~19_combout\,
	combout => \ShiftRight1~48_combout\);

-- Location: FF_X71_Y7_N44
\Selector22~0_OTERM475_NEW_REG746\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~48_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector22~0_OTERM475_OTERM747\);

-- Location: MLABCELL_X72_Y7_N27
\ShiftRight0~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight0~11_combout\ = ( \Mux223~0_combout\ & ( \Mux224~0_combout\ & ( (!\NxR.aluData2[1]~17_combout\ & (!\NxR.aluData2[3]~18_combout\ & \NxR.aluData2[2]~19_combout\)) ) ) ) # ( !\Mux223~0_combout\ & ( \Mux224~0_combout\ & ( 
-- (!\NxR.aluData2[0]~16_combout\ & (!\NxR.aluData2[1]~17_combout\ & (!\NxR.aluData2[3]~18_combout\ & \NxR.aluData2[2]~19_combout\))) ) ) ) # ( \Mux223~0_combout\ & ( !\Mux224~0_combout\ & ( (\NxR.aluData2[0]~16_combout\ & (!\NxR.aluData2[1]~17_combout\ & 
-- (!\NxR.aluData2[3]~18_combout\ & \NxR.aluData2[2]~19_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000100000000000000100000000000000011000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datab => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datac => \ALT_INV_NxR.aluData2[3]~18_combout\,
	datad => \ALT_INV_NxR.aluData2[2]~19_combout\,
	datae => \ALT_INV_Mux223~0_combout\,
	dataf => \ALT_INV_Mux224~0_combout\,
	combout => \ShiftRight0~11_combout\);

-- Location: FF_X72_Y7_N28
\Selector22~0_OTERM475_NEW_REG748\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight0~11_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector22~0_OTERM475_OTERM749\);

-- Location: LABCELL_X79_Y7_N30
\Selector22~0_RTM0477\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector22~0_RTM0477_combout\ = ( \R.aluOp.ALUOpSRA~q\ & ( \Selector22~0_OTERM475_OTERM749\ & ( (((\ShiftRight1~27_OTERM19\ & !\ShiftRight0~7_OTERM233DUPLICATE_q\)) # (\R.aluOp.ALUOpSRL~q\)) # (\Selector22~0_OTERM475_OTERM747\) ) ) ) # ( 
-- !\R.aluOp.ALUOpSRA~q\ & ( \Selector22~0_OTERM475_OTERM749\ & ( \R.aluOp.ALUOpSRL~q\ ) ) ) # ( \R.aluOp.ALUOpSRA~q\ & ( !\Selector22~0_OTERM475_OTERM749\ & ( ((\ShiftRight1~27_OTERM19\ & !\ShiftRight0~7_OTERM233DUPLICATE_q\)) # 
-- (\Selector22~0_OTERM475_OTERM747\) ) ) ) # ( !\R.aluOp.ALUOpSRA~q\ & ( !\Selector22~0_OTERM475_OTERM749\ & ( (\ShiftRight1~27_OTERM19\ & (\R.aluOp.ALUOpSRL~q\ & !\ShiftRight0~7_OTERM233DUPLICATE_q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000000011101110101010100001111000011110111111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector22~0_OTERM475_OTERM747\,
	datab => \ALT_INV_ShiftRight1~27_OTERM19\,
	datac => \ALT_INV_R.aluOp.ALUOpSRL~q\,
	datad => \ALT_INV_ShiftRight0~7_OTERM233DUPLICATE_q\,
	datae => \ALT_INV_R.aluOp.ALUOpSRA~q\,
	dataf => \ALT_INV_Selector22~0_OTERM475_OTERM749\,
	combout => \Selector22~0_RTM0477_combout\);

-- Location: MLABCELL_X78_Y7_N54
\ShiftLeft0~46\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~46_combout\ = ( \R.aluData2\(2) & ( \R.aluData2\(3) & ( \ShiftLeft0~20_OTERM291\ ) ) ) # ( !\R.aluData2\(2) & ( \R.aluData2\(3) & ( \ShiftLeft0~28_OTERM295\ ) ) ) # ( \R.aluData2\(2) & ( !\R.aluData2\(3) & ( \ShiftLeft0~36_OTERM603\ ) ) ) # ( 
-- !\R.aluData2\(2) & ( !\R.aluData2\(3) & ( \ShiftLeft0~45_OTERM757\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110011010101010101010100001111000011110000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~36_OTERM603\,
	datab => \ALT_INV_ShiftLeft0~45_OTERM757\,
	datac => \ALT_INV_ShiftLeft0~28_OTERM295\,
	datad => \ALT_INV_ShiftLeft0~20_OTERM291\,
	datae => \ALT_INV_R.aluData2\(2),
	dataf => \ALT_INV_R.aluData2\(3),
	combout => \ShiftLeft0~46_combout\);

-- Location: LABCELL_X77_Y8_N54
\Selector6~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector6~0_combout\ = ( \R.aluOp.ALUOpXor~DUPLICATE_q\ & ( !\Selector17~0_OTERM391\ & ( (!\R.aluData1\(26) & (((!\R.aluData2\(26))))) # (\R.aluData1\(26) & (!\R.aluOp.ALUOpAnd~DUPLICATE_q\ & (!\R.aluOp.ALUOpOr~q\ & \R.aluData2\(26)))) ) ) ) # ( 
-- !\R.aluOp.ALUOpXor~DUPLICATE_q\ & ( !\Selector17~0_OTERM391\ & ( (!\R.aluOp.ALUOpOr~q\ & ((!\R.aluOp.ALUOpAnd~DUPLICATE_q\) # ((!\R.aluData1\(26)) # (!\R.aluData2\(26))))) # (\R.aluOp.ALUOpOr~q\ & (((!\R.aluData1\(26) & !\R.aluData2\(26))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111110011001000111100000000100000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpAnd~DUPLICATE_q\,
	datab => \ALT_INV_R.aluOp.ALUOpOr~q\,
	datac => \ALT_INV_R.aluData1\(26),
	datad => \ALT_INV_R.aluData2\(26),
	datae => \ALT_INV_R.aluOp.ALUOpXor~DUPLICATE_q\,
	dataf => \ALT_INV_Selector17~0_OTERM391\,
	combout => \Selector6~0_combout\);

-- Location: MLABCELL_X78_Y7_N51
\ShiftLeft0~44\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~44_combout\ = ( \R.aluData2\(3) & ( (\ShiftLeft0~2_OTERM221\ & !\R.aluData2\(2)) ) ) # ( !\R.aluData2\(3) & ( (!\R.aluData2\(2) & ((\ShiftLeft0~13_OTERM285\))) # (\R.aluData2\(2) & (\ShiftLeft0~8_OTERM207\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001111001111000000111100111101000100010001000100010001000100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~2_OTERM221\,
	datab => \ALT_INV_R.aluData2\(2),
	datac => \ALT_INV_ShiftLeft0~8_OTERM207\,
	datad => \ALT_INV_ShiftLeft0~13_OTERM285\,
	dataf => \ALT_INV_R.aluData2\(3),
	combout => \ShiftLeft0~44_combout\);

-- Location: LABCELL_X77_Y7_N12
\Selector6~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector6~1_combout\ = ( \Selector6~0_combout\ & ( \ShiftLeft0~44_combout\ & ( (!\R.aluData2\(4) & (!\Selector22~0_RTM0477_combout\ & ((!\R.aluOp.ALUOpSLL~q\) # (!\ShiftLeft0~46_combout\)))) # (\R.aluData2\(4) & (((!\R.aluOp.ALUOpSLL~q\)))) ) ) ) # ( 
-- \Selector6~0_combout\ & ( !\ShiftLeft0~44_combout\ & ( ((!\Selector22~0_RTM0477_combout\ & ((!\R.aluOp.ALUOpSLL~q\) # (!\ShiftLeft0~46_combout\)))) # (\R.aluData2\(4)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101011111000111100000000000000001010110010001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector22~0_RTM0477_combout\,
	datab => \ALT_INV_R.aluOp.ALUOpSLL~q\,
	datac => \ALT_INV_R.aluData2\(4),
	datad => \ALT_INV_ShiftLeft0~46_combout\,
	datae => \ALT_INV_Selector6~0_combout\,
	dataf => \ALT_INV_ShiftLeft0~44_combout\,
	combout => \Selector6~1_combout\);

-- Location: MLABCELL_X78_Y7_N15
\Selector6~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector6~2_combout\ = ( \Add2~105_sumout\ & ( (!\Selector6~1_combout\) # (((\Add1~105_sumout\ & \R.aluOp.ALUOpAdd~q\)) # (\R.aluOp.ALUOpSub~q\)) ) ) # ( !\Add2~105_sumout\ & ( (!\Selector6~1_combout\) # ((\Add1~105_sumout\ & \R.aluOp.ALUOpAdd~q\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010101110101011101010111010101110101011111111111010101111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector6~1_combout\,
	datab => \ALT_INV_Add1~105_sumout\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_R.aluOp.ALUOpSub~q\,
	dataf => \ALT_INV_Add2~105_sumout\,
	combout => \Selector6~2_combout\);

-- Location: FF_X78_Y7_N17
\R.aluRes[26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector6~2_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(26));

-- Location: MLABCELL_X78_Y7_N48
\vAluRes~28\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~28_combout\ = ( \R.aluRes\(26) & ( !\R.aluCalc~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011110000111100001111000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_R.aluCalc~q\,
	dataf => \ALT_INV_R.aluRes\(26),
	combout => \vAluRes~28_combout\);

-- Location: MLABCELL_X78_Y7_N24
\Comb:vJumpAdr[26]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[26]~0_combout\ = ( \Add3~105_sumout\ & ( (!\Equal4~2_combout\) # ((\vAluRes~27_combout\) # (\vAluRes~28_combout\)) ) ) # ( !\Add3~105_sumout\ & ( (\Equal4~2_combout\ & ((\vAluRes~27_combout\) # (\vAluRes~28_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010101010101000001010101010110101111111111111010111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Equal4~2_combout\,
	datac => \ALT_INV_vAluRes~28_combout\,
	datad => \ALT_INV_vAluRes~27_combout\,
	dataf => \ALT_INV_Add3~105_sumout\,
	combout => \Comb:vJumpAdr[26]~0_combout\);

-- Location: FF_X78_Y7_N25
\R.curPC[26]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[26]~0_combout\,
	asdata => \Add0~97_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(26));

-- Location: LABCELL_X81_Y5_N45
\Add0~101\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add0~101_sumout\ = SUM(( \R.curPC\(27) ) + ( GND ) + ( \Add0~98\ ))
-- \Add0~102\ = CARRY(( \R.curPC\(27) ) + ( GND ) + ( \Add0~98\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curPC\(27),
	cin => \Add0~98\,
	sumout => \Add0~101_sumout\,
	cout => \Add0~102\);

-- Location: IOIBUF_X84_Y0_N52
\avm_d_readdata[3]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(3),
	o => \avm_d_readdata[3]~input_o\);

-- Location: LABCELL_X81_Y5_N24
\Comb:vRegWriteData[27]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[27]~1_combout\ = ( \Add1~109_sumout\ & ( \R.curInst\(13) & ( (!\R.memToReg~q\ & (((\R.aluOp.ALUOpAdd~q\)))) # (\R.memToReg~q\ & (!\R.curInst\(14) & ((\avm_d_readdata[3]~input_o\)))) ) ) ) # ( !\Add1~109_sumout\ & ( \R.curInst\(13) & ( 
-- (!\R.curInst\(14) & (\R.memToReg~q\ & \avm_d_readdata[3]~input_o\)) ) ) ) # ( \Add1~109_sumout\ & ( !\R.curInst\(13) & ( (!\R.memToReg~q\ & ((\R.aluOp.ALUOpAdd~q\))) # (\R.memToReg~q\ & (!\R.curInst\(14))) ) ) ) # ( !\Add1~109_sumout\ & ( !\R.curInst\(13) 
-- & ( (!\R.curInst\(14) & \R.memToReg~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010001000100010001011100010111000000000001000100000110000101110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(14),
	datab => \ALT_INV_R.memToReg~q\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_avm_d_readdata[3]~input_o\,
	datae => \ALT_INV_Add1~109_sumout\,
	dataf => \ALT_INV_R.curInst\(13),
	combout => \Comb:vRegWriteData[27]~1_combout\);

-- Location: FF_X79_Y4_N13
\R.aluRes[27]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector5~5_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes[27]~DUPLICATE_q\);

-- Location: LABCELL_X80_Y4_N30
\Comb:vRegWriteData[27]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[27]~3_combout\ = ( \Selector5~2_combout\ & ( (!\R.aluRes[27]~DUPLICATE_q\ & (!\R.aluCalc~q\ & !\R.memToReg~q\)) ) ) # ( !\Selector5~2_combout\ & ( (!\R.aluCalc~q\ & (!\R.aluRes[27]~DUPLICATE_q\ & (!\R.memToReg~q\))) # (\R.aluCalc~q\ & 
-- (((\Selector5~4_combout\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000000010110011100000001011001110000000100000001000000010000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluRes[27]~DUPLICATE_q\,
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_R.memToReg~q\,
	datad => \ALT_INV_Selector5~4_combout\,
	dataf => \ALT_INV_Selector5~2_combout\,
	combout => \Comb:vRegWriteData[27]~3_combout\);

-- Location: LABCELL_X79_Y1_N24
\Comb:vRegWriteData[27]~2_RESYN1108\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[27]~2_RESYN1108_BDD1109\ = ( \R.curInst\(12) & ( !\avm_d_readdata[23]~input_o\ ) ) # ( !\R.curInst\(12) & ( !\avm_d_readdata[31]~input_o\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1100110011001100110011001100110011110000111100001111000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_avm_d_readdata[31]~input_o\,
	datac => \ALT_INV_avm_d_readdata[23]~input_o\,
	dataf => \ALT_INV_R.curInst\(12),
	combout => \Comb:vRegWriteData[27]~2_RESYN1108_BDD1109\);

-- Location: LABCELL_X79_Y1_N45
\Comb:vRegWriteData[27]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[27]~2_combout\ = ( \avm_d_readdata[3]~input_o\ & ( \Comb:vRegWriteData[27]~2_RESYN1108_BDD1109\ & ( (\R.memToReg~q\ & (((!\R.curInst\(13)) # (\R.curInst\(12))) # (\R.curInst\(14)))) ) ) ) # ( !\avm_d_readdata[3]~input_o\ & ( 
-- \Comb:vRegWriteData[27]~2_RESYN1108_BDD1109\ & ( \R.memToReg~q\ ) ) ) # ( \avm_d_readdata[3]~input_o\ & ( !\Comb:vRegWriteData[27]~2_RESYN1108_BDD1109\ & ( (\R.memToReg~q\ & (((\R.curInst\(13) & \R.curInst\(12))) # (\R.curInst\(14)))) ) ) ) # ( 
-- !\avm_d_readdata[3]~input_o\ & ( !\Comb:vRegWriteData[27]~2_RESYN1108_BDD1109\ & ( (\R.memToReg~q\ & ((\R.curInst\(13)) # (\R.curInst\(14)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000011100000111000001010000011100001111000011110000110100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(14),
	datab => \ALT_INV_R.curInst\(13),
	datac => \ALT_INV_R.memToReg~q\,
	datad => \ALT_INV_R.curInst\(12),
	datae => \ALT_INV_avm_d_readdata[3]~input_o\,
	dataf => \ALT_INV_Comb:vRegWriteData[27]~2_RESYN1108_BDD1109\,
	combout => \Comb:vRegWriteData[27]~2_combout\);

-- Location: LABCELL_X81_Y5_N6
\Comb:vRegWriteData[27]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[27]~0_combout\ = ( \Comb:vRegWriteData[27]~3_combout\ & ( !\Comb:vRegWriteData[27]~2_combout\ & ( (\R.aluCalc~q\ & (((\Add2~109_sumout\ & \R.aluOp.ALUOpSub~q\)) # (\Comb:vRegWriteData[27]~1_combout\))) ) ) ) # ( 
-- !\Comb:vRegWriteData[27]~3_combout\ & ( !\Comb:vRegWriteData[27]~2_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111000000000001111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add2~109_sumout\,
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_Comb:vRegWriteData[27]~1_combout\,
	datad => \ALT_INV_R.aluCalc~q\,
	datae => \ALT_INV_Comb:vRegWriteData[27]~3_combout\,
	dataf => \ALT_INV_Comb:vRegWriteData[27]~2_combout\,
	combout => \Comb:vRegWriteData[27]~0_combout\);

-- Location: FF_X81_Y5_N47
\R.regWriteData[27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Add0~101_sumout\,
	asdata => \Comb:vRegWriteData[27]~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(27));

-- Location: FF_X71_Y4_N26
\RegFile[29][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(27),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][27]~q\);

-- Location: FF_X67_Y4_N55
\RegFile[26][27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[26][27]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][27]~q\);

-- Location: LABCELL_X71_Y4_N48
\Mux95~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux95~22_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[24][27]~q\))) # (\R.curInst\(20) & (\RegFile[25][27]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & (\RegFile[26][27]~q\)) # (\R.curInst\(20) & ((\RegFile[27][27]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[25][27]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[26][27]~q\,
	datad => \ALT_INV_RegFile[27][27]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][27]~q\,
	combout => \Mux95~22_combout\);

-- Location: LABCELL_X71_Y4_N24
\Mux95~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux95~9_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux95~22_combout\)))) # (\R.curInst\(22) & ((!\Mux95~22_combout\ & ((\RegFile[28][27]~q\))) # (\Mux95~22_combout\ & (\RegFile[29][27]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux95~22_combout\)))) # (\R.curInst\(22) & ((!\Mux95~22_combout\ & ((\RegFile[30][27]~q\))) # (\Mux95~22_combout\ & (\RegFile[31][27]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[29][27]~q\,
	datab => \ALT_INV_RegFile[31][27]~q\,
	datac => \ALT_INV_RegFile[30][27]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux95~22_combout\,
	datag => \ALT_INV_RegFile[28][27]~q\,
	combout => \Mux95~9_combout\);

-- Location: MLABCELL_X65_Y6_N18
\Mux95~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux95~0_combout\ = ( \RegFile[6][27]~q\ & ( \R.curInst\(20) & ( (!\R.curInst\(21) & ((\RegFile[5][27]~q\))) # (\R.curInst\(21) & (\RegFile[7][27]~q\)) ) ) ) # ( !\RegFile[6][27]~q\ & ( \R.curInst\(20) & ( (!\R.curInst\(21) & ((\RegFile[5][27]~q\))) # 
-- (\R.curInst\(21) & (\RegFile[7][27]~q\)) ) ) ) # ( \RegFile[6][27]~q\ & ( !\R.curInst\(20) & ( (\R.curInst\(21)) # (\RegFile[4][27]~q\) ) ) ) # ( !\RegFile[6][27]~q\ & ( !\R.curInst\(20) & ( (\RegFile[4][27]~q\ & !\R.curInst\(21)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100010001000100011101110111011100000011110011110000001111001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[4][27]~q\,
	datab => \ALT_INV_R.curInst\(21),
	datac => \ALT_INV_RegFile[7][27]~q\,
	datad => \ALT_INV_RegFile[5][27]~q\,
	datae => \ALT_INV_RegFile[6][27]~q\,
	dataf => \ALT_INV_R.curInst\(20),
	combout => \Mux95~0_combout\);

-- Location: LABCELL_X66_Y4_N42
\Mux95~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux95~26_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (\R.curInst\(20) & (\RegFile[1][27]~q\))) # (\R.curInst\(22) & (((\Mux95~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (((\RegFile[2][27]~q\)))) # 
-- (\R.curInst\(20) & (\RegFile[3][27]~q\)))) # (\R.curInst\(22) & ((((\Mux95~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000000000111010000000000000011111111110001110111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][27]~q\,
	datab => \ALT_INV_R.curInst\(20),
	datac => \ALT_INV_RegFile[2][27]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux95~0_combout\,
	datag => \ALT_INV_RegFile[1][27]~q\,
	combout => \Mux95~26_combout\);

-- Location: LABCELL_X66_Y4_N6
\Mux95~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux95~18_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & (\RegFile[16][27]~q\)) # (\R.curInst\(20) & ((\RegFile[17][27]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & ((\RegFile[18][27]~q\))) # (\R.curInst\(20) & (\RegFile[19][27]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110000110011111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[19][27]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[18][27]~q\,
	datad => \ALT_INV_RegFile[17][27]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][27]~q\,
	combout => \Mux95~18_combout\);

-- Location: LABCELL_X70_Y4_N24
\Mux95~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux95~5_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux95~18_combout\))))) # (\R.curInst\(22) & (((!\Mux95~18_combout\ & ((\RegFile[20][27]~q\))) # (\Mux95~18_combout\ & (\RegFile[21][27]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux95~18_combout\)))) # (\R.curInst\(22) & ((!\Mux95~18_combout\ & (\RegFile[22][27]~q\)) # (\Mux95~18_combout\ & ((\RegFile[23][27]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][27]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[22][27]~q\,
	datad => \ALT_INV_RegFile[23][27]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux95~18_combout\,
	datag => \ALT_INV_RegFile[20][27]~q\,
	combout => \Mux95~5_combout\);

-- Location: LABCELL_X67_Y8_N0
\Mux95~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux95~14_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[8][27]~q\))) # (\R.curInst\(20) & (\RegFile[9][27]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & (\RegFile[10][27]~q\)) # (\R.curInst\(20) & ((\RegFile[11][27]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][27]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[10][27]~q\,
	datad => \ALT_INV_RegFile[11][27]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][27]~q\,
	combout => \Mux95~14_combout\);

-- Location: LABCELL_X71_Y4_N54
\Mux95~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux95~1_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux95~14_combout\))))) # (\R.curInst\(22) & (((!\Mux95~14_combout\ & ((\RegFile[12][27]~q\))) # (\Mux95~14_combout\ & (\RegFile[13][27]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux95~14_combout\)))) # (\R.curInst\(22) & ((!\Mux95~14_combout\ & (\RegFile[14][27]~q\)) # (\Mux95~14_combout\ & ((\RegFile[15][27]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][27]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[14][27]~q\,
	datad => \ALT_INV_RegFile[15][27]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux95~14_combout\,
	datag => \ALT_INV_RegFile[12][27]~q\,
	combout => \Mux95~1_combout\);

-- Location: MLABCELL_X72_Y4_N45
\Mux95~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux95~13_combout\ = ( \Mux95~5_combout\ & ( \Mux95~1_combout\ & ( (!\R.curInst\(24) & (((\Mux95~26_combout\)) # (\R.curInst\(23)))) # (\R.curInst\(24) & ((!\R.curInst\(23)) # ((\Mux95~9_combout\)))) ) ) ) # ( !\Mux95~5_combout\ & ( \Mux95~1_combout\ & ( 
-- (!\R.curInst\(24) & (((\Mux95~26_combout\)) # (\R.curInst\(23)))) # (\R.curInst\(24) & (\R.curInst\(23) & (\Mux95~9_combout\))) ) ) ) # ( \Mux95~5_combout\ & ( !\Mux95~1_combout\ & ( (!\R.curInst\(24) & (!\R.curInst\(23) & ((\Mux95~26_combout\)))) # 
-- (\R.curInst\(24) & ((!\R.curInst\(23)) # ((\Mux95~9_combout\)))) ) ) ) # ( !\Mux95~5_combout\ & ( !\Mux95~1_combout\ & ( (!\R.curInst\(24) & (!\R.curInst\(23) & ((\Mux95~26_combout\)))) # (\R.curInst\(24) & (\R.curInst\(23) & (\Mux95~9_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000110001001010001011100110100100011101010110110011111101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(24),
	datab => \ALT_INV_R.curInst\(23),
	datac => \ALT_INV_Mux95~9_combout\,
	datad => \ALT_INV_Mux95~26_combout\,
	datae => \ALT_INV_Mux95~5_combout\,
	dataf => \ALT_INV_Mux95~1_combout\,
	combout => \Mux95~13_combout\);

-- Location: LABCELL_X73_Y4_N0
\NxR.aluData2[27]~24\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[27]~24_combout\ = ( \Mux95~13_combout\ & ( (!\vAluSrc2~1_combout\) # ((\Equal4~1_combout\ & \Mux127~0_combout\)) ) ) # ( !\Mux95~13_combout\ & ( (\vAluSrc2~1_combout\ & (\Equal4~1_combout\ & \Mux127~0_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000100000001000000010000000110101011101010111010101110101011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluSrc2~1_combout\,
	datab => \ALT_INV_Equal4~1_combout\,
	datac => \ALT_INV_Mux127~0_combout\,
	dataf => \ALT_INV_Mux95~13_combout\,
	combout => \NxR.aluData2[27]~24_combout\);

-- Location: FF_X73_Y4_N22
\R.aluData2[27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \NxR.aluData2[27]~24_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData2\(27));

-- Location: LABCELL_X79_Y5_N42
\Comb:vJumpAdr[27]~0_RESYN1030\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[27]~0_RESYN1030_BDD1031\ = ( \R.aluRes[27]~DUPLICATE_q\ & ( \Selector5~2_combout\ ) ) # ( !\R.aluRes[27]~DUPLICATE_q\ & ( \Selector5~2_combout\ & ( \R.aluCalc~q\ ) ) ) # ( \R.aluRes[27]~DUPLICATE_q\ & ( !\Selector5~2_combout\ & ( 
-- (!\R.aluCalc~q\) # ((!\Selector5~4_combout\) # ((\Add2~109_sumout\ & \R.aluOp.ALUOpSub~q\))) ) ) ) # ( !\R.aluRes[27]~DUPLICATE_q\ & ( !\Selector5~2_combout\ & ( (\R.aluCalc~q\ & ((!\Selector5~4_combout\) # ((\Add2~109_sumout\ & \R.aluOp.ALUOpSub~q\)))) ) 
-- ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100010001000101111011101110111101010101010101011111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluCalc~q\,
	datab => \ALT_INV_Selector5~4_combout\,
	datac => \ALT_INV_Add2~109_sumout\,
	datad => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datae => \ALT_INV_R.aluRes[27]~DUPLICATE_q\,
	dataf => \ALT_INV_Selector5~2_combout\,
	combout => \Comb:vJumpAdr[27]~0_RESYN1030_BDD1031\);

-- Location: LABCELL_X80_Y4_N12
\Comb:vJumpAdr[27]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[27]~0_combout\ = ( \Equal4~2_combout\ & ( \Add3~109_sumout\ & ( ((\Add1~109_sumout\ & (\R.aluOp.ALUOpAdd~q\ & \R.aluCalc~q\))) # (\Comb:vJumpAdr[27]~0_RESYN1030_BDD1031\) ) ) ) # ( !\Equal4~2_combout\ & ( \Add3~109_sumout\ ) ) # ( 
-- \Equal4~2_combout\ & ( !\Add3~109_sumout\ & ( ((\Add1~109_sumout\ & (\R.aluOp.ALUOpAdd~q\ & \R.aluCalc~q\))) # (\Comb:vJumpAdr[27]~0_RESYN1030_BDD1031\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110001111111111111111111110000111100011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add1~109_sumout\,
	datab => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datac => \ALT_INV_Comb:vJumpAdr[27]~0_RESYN1030_BDD1031\,
	datad => \ALT_INV_R.aluCalc~q\,
	datae => \ALT_INV_Equal4~2_combout\,
	dataf => \ALT_INV_Add3~109_sumout\,
	combout => \Comb:vJumpAdr[27]~0_combout\);

-- Location: FF_X80_Y4_N13
\R.curPC[27]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[27]~0_combout\,
	asdata => \Add0~101_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(27));

-- Location: IOIBUF_X34_Y0_N75
\avm_d_readdata[4]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(4),
	o => \avm_d_readdata[4]~input_o\);

-- Location: LABCELL_X79_Y2_N36
\Comb:vRegWriteData[28]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[28]~1_combout\ = ( \avm_d_readdata[23]~input_o\ & ( \avm_d_readdata[4]~input_o\ & ( (!\R.curInst\(14) & ((!\R.curInst\(12) & ((\avm_d_readdata[31]~input_o\) # (\R.curInst\(13)))) # (\R.curInst\(12) & (!\R.curInst\(13))))) ) ) ) # ( 
-- !\avm_d_readdata[23]~input_o\ & ( \avm_d_readdata[4]~input_o\ & ( (!\R.curInst\(12) & (!\R.curInst\(14) & ((\avm_d_readdata[31]~input_o\) # (\R.curInst\(13))))) ) ) ) # ( \avm_d_readdata[23]~input_o\ & ( !\avm_d_readdata[4]~input_o\ & ( (!\R.curInst\(14) 
-- & (!\R.curInst\(13) & ((\avm_d_readdata[31]~input_o\) # (\R.curInst\(12))))) ) ) ) # ( !\avm_d_readdata[23]~input_o\ & ( !\avm_d_readdata[4]~input_o\ & ( (!\R.curInst\(12) & (!\R.curInst\(14) & (!\R.curInst\(13) & \avm_d_readdata[31]~input_o\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000010000000010000001100000000001000100010000100100011001000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(12),
	datab => \ALT_INV_R.curInst\(14),
	datac => \ALT_INV_R.curInst\(13),
	datad => \ALT_INV_avm_d_readdata[31]~input_o\,
	datae => \ALT_INV_avm_d_readdata[23]~input_o\,
	dataf => \ALT_INV_avm_d_readdata[4]~input_o\,
	combout => \Comb:vRegWriteData[28]~1_combout\);

-- Location: MLABCELL_X78_Y4_N30
\Comb:vRegWriteData[28]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[28]~2_combout\ = ( \Comb:vRegWriteData[28]~1_combout\ & ( (!\Selector4~1_combout\ & (!\R.memToReg~q\ & ((!\R.aluOp.ALUOpAdd~q\) # (!\Add1~113_sumout\)))) ) ) # ( !\Comb:vRegWriteData[28]~1_combout\ & ( ((!\Selector4~1_combout\ & 
-- ((!\R.aluOp.ALUOpAdd~q\) # (!\Add1~113_sumout\)))) # (\R.memToReg~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1100111110001111110011111000111111000000100000001100000010000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datab => \ALT_INV_Selector4~1_combout\,
	datac => \ALT_INV_R.memToReg~q\,
	datad => \ALT_INV_Add1~113_sumout\,
	dataf => \ALT_INV_Comb:vRegWriteData[28]~1_combout\,
	combout => \Comb:vRegWriteData[28]~2_combout\);

-- Location: MLABCELL_X78_Y4_N18
\Comb:vRegWriteData[28]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[28]~0_combout\ = ( \R.memToReg~q\ & ( \Add2~113_sumout\ & ( !\Comb:vRegWriteData[28]~2_combout\ ) ) ) # ( !\R.memToReg~q\ & ( \Add2~113_sumout\ & ( (!\R.aluCalc~q\ & (((\R.aluRes\(28))))) # (\R.aluCalc~q\ & 
-- (((!\Comb:vRegWriteData[28]~2_combout\)) # (\R.aluOp.ALUOpSub~q\))) ) ) ) # ( \R.memToReg~q\ & ( !\Add2~113_sumout\ & ( !\Comb:vRegWriteData[28]~2_combout\ ) ) ) # ( !\R.memToReg~q\ & ( !\Add2~113_sumout\ & ( (!\R.aluCalc~q\ & (\R.aluRes\(28))) # 
-- (\R.aluCalc~q\ & ((!\Comb:vRegWriteData[28]~2_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101111100001010111111110000000001011111000110111111111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluCalc~q\,
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_R.aluRes\(28),
	datad => \ALT_INV_Comb:vRegWriteData[28]~2_combout\,
	datae => \ALT_INV_R.memToReg~q\,
	dataf => \ALT_INV_Add2~113_sumout\,
	combout => \Comb:vRegWriteData[28]~0_combout\);

-- Location: FF_X81_Y5_N50
\R.regWriteData[28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Add0~105_sumout\,
	asdata => \Comb:vRegWriteData[28]~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(28));

-- Location: FF_X65_Y1_N38
\RegFile[13][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(28),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~7_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[13][28]~q\);

-- Location: FF_X65_Y1_N14
\RegFile[15][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(28),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][28]~q\);

-- Location: LABCELL_X55_Y1_N12
\RegFile[14][28]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[14][28]~feeder_combout\ = ( \R.regWriteData\(28) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(28),
	combout => \RegFile[14][28]~feeder_combout\);

-- Location: FF_X55_Y1_N13
\RegFile[14][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[14][28]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][28]~q\);

-- Location: FF_X65_Y1_N50
\RegFile[11][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(28),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~20_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[11][28]~q\);

-- Location: LABCELL_X71_Y8_N21
\RegFile[9][28]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[9][28]~feeder_combout\ = ( \R.regWriteData\(28) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(28),
	combout => \RegFile[9][28]~feeder_combout\);

-- Location: FF_X71_Y8_N22
\RegFile[9][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[9][28]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~19_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[9][28]~q\);

-- Location: LABCELL_X57_Y1_N30
\RegFile[10][28]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[10][28]~feeder_combout\ = ( \R.regWriteData\(28) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(28),
	combout => \RegFile[10][28]~feeder_combout\);

-- Location: FF_X57_Y1_N31
\RegFile[10][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[10][28]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~22_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[10][28]~q\);

-- Location: MLABCELL_X59_Y1_N12
\RegFile[8][28]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[8][28]~feeder_combout\ = ( \R.regWriteData\(28) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(28),
	combout => \RegFile[8][28]~feeder_combout\);

-- Location: FF_X59_Y1_N14
\RegFile[8][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[8][28]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~21_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[8][28]~q\);

-- Location: MLABCELL_X65_Y1_N24
\Mux94~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux94~14_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[8][28]~q\))) # (\R.curInst\(20) & (\RegFile[9][28]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[10][28]~q\))) # (\R.curInst\(20) & (\RegFile[11][28]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[11][28]~q\,
	datab => \ALT_INV_RegFile[9][28]~q\,
	datac => \ALT_INV_RegFile[10][28]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][28]~q\,
	combout => \Mux94~14_combout\);

-- Location: LABCELL_X57_Y1_N9
\RegFile[12][28]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[12][28]~feeder_combout\ = ( \R.regWriteData\(28) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(28),
	combout => \RegFile[12][28]~feeder_combout\);

-- Location: FF_X57_Y1_N10
\RegFile[12][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[12][28]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][28]~q\);

-- Location: MLABCELL_X65_Y1_N12
\Mux94~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux94~1_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux94~14_combout\)))) # (\R.curInst\(22) & ((!\Mux94~14_combout\ & ((\RegFile[12][28]~q\))) # (\Mux94~14_combout\ & (\RegFile[13][28]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux94~14_combout\)))) # (\R.curInst\(22) & ((!\Mux94~14_combout\ & ((\RegFile[14][28]~q\))) # (\Mux94~14_combout\ & (\RegFile[15][28]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][28]~q\,
	datab => \ALT_INV_RegFile[15][28]~q\,
	datac => \ALT_INV_RegFile[14][28]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux94~14_combout\,
	datag => \ALT_INV_RegFile[12][28]~q\,
	combout => \Mux94~1_combout\);

-- Location: FF_X71_Y5_N19
\RegFile[31][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(28),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][28]~q\);

-- Location: FF_X68_Y6_N1
\RegFile[29][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(28),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~15_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[29][28]~q\);

-- Location: FF_X57_Y6_N13
\RegFile[30][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(28),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~18_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[30][28]~q\);

-- Location: FF_X67_Y4_N20
\RegFile[27][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(28),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~28_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[27][28]~q\);

-- Location: FF_X67_Y4_N26
\RegFile[25][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(28),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~27_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[25][28]~q\);

-- Location: LABCELL_X67_Y4_N48
\RegFile[26][28]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[26][28]~feeder_combout\ = ( \R.regWriteData\(28) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(28),
	combout => \RegFile[26][28]~feeder_combout\);

-- Location: FF_X67_Y4_N50
\RegFile[26][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[26][28]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~30_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[26][28]~q\);

-- Location: LABCELL_X56_Y2_N15
\RegFile[24][28]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[24][28]~feeder_combout\ = ( \R.regWriteData\(28) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(28),
	combout => \RegFile[24][28]~feeder_combout\);

-- Location: FF_X56_Y2_N16
\RegFile[24][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[24][28]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~29_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[24][28]~q\);

-- Location: LABCELL_X67_Y4_N24
\Mux94~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux94~22_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[24][28]~q\))) # (\R.curInst\(20) & (\RegFile[25][28]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[26][28]~q\))) # (\R.curInst\(20) & (\RegFile[27][28]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[27][28]~q\,
	datab => \ALT_INV_RegFile[25][28]~q\,
	datac => \ALT_INV_RegFile[26][28]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][28]~q\,
	combout => \Mux94~22_combout\);

-- Location: LABCELL_X71_Y8_N24
\RegFile[28][28]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[28][28]~feeder_combout\ = ( \R.regWriteData\(28) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(28),
	combout => \RegFile[28][28]~feeder_combout\);

-- Location: FF_X71_Y8_N25
\RegFile[28][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[28][28]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][28]~q\);

-- Location: LABCELL_X68_Y4_N12
\Mux94~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux94~9_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux94~22_combout\)))) # (\R.curInst\(22) & ((!\Mux94~22_combout\ & ((\RegFile[28][28]~q\))) # (\Mux94~22_combout\ & (\RegFile[29][28]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux94~22_combout\)))) # (\R.curInst\(22) & ((!\Mux94~22_combout\ & ((\RegFile[30][28]~q\))) # (\Mux94~22_combout\ & (\RegFile[31][28]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][28]~q\,
	datab => \ALT_INV_RegFile[29][28]~q\,
	datac => \ALT_INV_RegFile[30][28]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux94~22_combout\,
	datag => \ALT_INV_RegFile[28][28]~q\,
	combout => \Mux94~9_combout\);

-- Location: FF_X68_Y4_N2
\RegFile[3][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(28),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][28]~q\);

-- Location: FF_X71_Y5_N13
\RegFile[2][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(28),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][28]~q\);

-- Location: FF_X66_Y5_N1
\RegFile[5][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(28),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~1_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[5][28]~q\);

-- Location: LABCELL_X67_Y5_N21
\RegFile[4][28]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[4][28]~feeder_combout\ = ( \R.regWriteData\(28) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(28),
	combout => \RegFile[4][28]~feeder_combout\);

-- Location: FF_X67_Y5_N22
\RegFile[4][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[4][28]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[4][28]~q\);

-- Location: FF_X61_Y1_N38
\RegFile[7][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(28),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~3_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[7][28]~q\);

-- Location: FF_X61_Y1_N43
\RegFile[6][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(28),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][28]~q\);

-- Location: LABCELL_X67_Y4_N9
\Mux94~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux94~0_combout\ = ( \R.curInst\(21) & ( \R.curInst\(20) & ( \RegFile[7][28]~q\ ) ) ) # ( !\R.curInst\(21) & ( \R.curInst\(20) & ( \RegFile[5][28]~q\ ) ) ) # ( \R.curInst\(21) & ( !\R.curInst\(20) & ( \RegFile[6][28]~q\ ) ) ) # ( !\R.curInst\(21) & ( 
-- !\R.curInst\(20) & ( \RegFile[4][28]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110011000000001111111101010101010101010000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[5][28]~q\,
	datab => \ALT_INV_RegFile[4][28]~q\,
	datac => \ALT_INV_RegFile[7][28]~q\,
	datad => \ALT_INV_RegFile[6][28]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	combout => \Mux94~0_combout\);

-- Location: LABCELL_X71_Y8_N57
\RegFile[1][28]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[1][28]~feeder_combout\ = ( \R.regWriteData\(28) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(28),
	combout => \RegFile[1][28]~feeder_combout\);

-- Location: FF_X71_Y8_N59
\RegFile[1][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[1][28]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~5_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[1][28]~q\);

-- Location: LABCELL_X68_Y4_N0
\Mux94~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux94~26_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (\R.curInst\(20) & (\RegFile[1][28]~q\))) # (\R.curInst\(22) & (((\Mux94~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (((\RegFile[2][28]~q\)))) # 
-- (\R.curInst\(20) & (\RegFile[3][28]~q\)))) # (\R.curInst\(22) & ((((\Mux94~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000000000111010000000000000011111111110001110111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][28]~q\,
	datab => \ALT_INV_R.curInst\(20),
	datac => \ALT_INV_RegFile[2][28]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux94~0_combout\,
	datag => \ALT_INV_RegFile[1][28]~q\,
	combout => \Mux94~26_combout\);

-- Location: FF_X71_Y5_N37
\RegFile[23][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(28),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][28]~q\);

-- Location: LABCELL_X67_Y9_N54
\RegFile[21][28]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[21][28]~feeder_combout\ = ( \R.regWriteData\(28) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(28),
	combout => \RegFile[21][28]~feeder_combout\);

-- Location: FF_X67_Y9_N55
\RegFile[21][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[21][28]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~11_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[21][28]~q\);

-- Location: FF_X75_Y8_N43
\RegFile[22][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(28),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~14_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[22][28]~q\);

-- Location: FF_X67_Y9_N50
\RegFile[19][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(28),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~24_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[19][28]~q\);

-- Location: LABCELL_X67_Y9_N12
\RegFile[17][28]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[17][28]~feeder_combout\ = ( \R.regWriteData\(28) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(28),
	combout => \RegFile[17][28]~feeder_combout\);

-- Location: FF_X67_Y9_N14
\RegFile[17][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[17][28]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~23_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[17][28]~q\);

-- Location: LABCELL_X63_Y10_N15
\RegFile[18][28]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[18][28]~feeder_combout\ = ( \R.regWriteData\(28) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(28),
	combout => \RegFile[18][28]~feeder_combout\);

-- Location: FF_X63_Y10_N16
\RegFile[18][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][28]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][28]~q\);

-- Location: LABCELL_X63_Y9_N21
\RegFile[16][28]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[16][28]~feeder_combout\ = ( \R.regWriteData\(28) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(28),
	combout => \RegFile[16][28]~feeder_combout\);

-- Location: FF_X63_Y9_N22
\RegFile[16][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[16][28]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][28]~q\);

-- Location: LABCELL_X67_Y6_N33
\Mux94~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux94~18_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[16][28]~q\))) # (\R.curInst\(20) & (\RegFile[17][28]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[18][28]~q\))) # (\R.curInst\(20) & (\RegFile[19][28]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[19][28]~q\,
	datab => \ALT_INV_RegFile[17][28]~q\,
	datac => \ALT_INV_RegFile[18][28]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][28]~q\,
	combout => \Mux94~18_combout\);

-- Location: FF_X68_Y6_N34
\RegFile[20][28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(28),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~13_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[20][28]~q\);

-- Location: LABCELL_X67_Y6_N36
\Mux94~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux94~5_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux94~18_combout\)))) # (\R.curInst\(22) & ((!\Mux94~18_combout\ & ((\RegFile[20][28]~q\))) # (\Mux94~18_combout\ & (\RegFile[21][28]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux94~18_combout\)))) # (\R.curInst\(22) & ((!\Mux94~18_combout\ & ((\RegFile[22][28]~q\))) # (\Mux94~18_combout\ & (\RegFile[23][28]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[23][28]~q\,
	datab => \ALT_INV_RegFile[21][28]~q\,
	datac => \ALT_INV_RegFile[22][28]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux94~18_combout\,
	datag => \ALT_INV_RegFile[20][28]~q\,
	combout => \Mux94~5_combout\);

-- Location: LABCELL_X68_Y4_N54
\Mux94~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux94~13_combout\ = ( \Mux94~26_combout\ & ( \Mux94~5_combout\ & ( (!\R.curInst\(23)) # ((!\R.curInst\(24) & (\Mux94~1_combout\)) # (\R.curInst\(24) & ((\Mux94~9_combout\)))) ) ) ) # ( !\Mux94~26_combout\ & ( \Mux94~5_combout\ & ( (!\R.curInst\(24) & 
-- (\R.curInst\(23) & (\Mux94~1_combout\))) # (\R.curInst\(24) & ((!\R.curInst\(23)) # ((\Mux94~9_combout\)))) ) ) ) # ( \Mux94~26_combout\ & ( !\Mux94~5_combout\ & ( (!\R.curInst\(24) & ((!\R.curInst\(23)) # ((\Mux94~1_combout\)))) # (\R.curInst\(24) & 
-- (\R.curInst\(23) & ((\Mux94~9_combout\)))) ) ) ) # ( !\Mux94~26_combout\ & ( !\Mux94~5_combout\ & ( (\R.curInst\(23) & ((!\R.curInst\(24) & (\Mux94~1_combout\)) # (\R.curInst\(24) & ((\Mux94~9_combout\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001000010011100010101001101101000110010101111100111011011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(24),
	datab => \ALT_INV_R.curInst\(23),
	datac => \ALT_INV_Mux94~1_combout\,
	datad => \ALT_INV_Mux94~9_combout\,
	datae => \ALT_INV_Mux94~26_combout\,
	dataf => \ALT_INV_Mux94~5_combout\,
	combout => \Mux94~13_combout\);

-- Location: LABCELL_X74_Y4_N54
\NxR.aluData2[28]~23\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[28]~23_combout\ = ( \Mux126~0_combout\ & ( (!\vAluSrc2~1_combout\ & ((\Mux94~13_combout\))) # (\vAluSrc2~1_combout\ & (\Equal4~1_combout\)) ) ) # ( !\Mux126~0_combout\ & ( (!\vAluSrc2~1_combout\ & \Mux94~13_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011110000000000001111000000000011111100110000001111110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Equal4~1_combout\,
	datac => \ALT_INV_vAluSrc2~1_combout\,
	datad => \ALT_INV_Mux94~13_combout\,
	dataf => \ALT_INV_Mux126~0_combout\,
	combout => \NxR.aluData2[28]~23_combout\);

-- Location: FF_X74_Y4_N56
\R.aluData2[28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR.aluData2[28]~23_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData2\(28));

-- Location: MLABCELL_X78_Y4_N48
\Comb:vJumpAdr[28]~0_RESYN1032\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[28]~0_RESYN1032_BDD1033\ = ( \Add2~113_sumout\ & ( ((\Add1~113_sumout\ & \R.aluOp.ALUOpAdd~q\)) # (\R.aluOp.ALUOpSub~q\) ) ) # ( !\Add2~113_sumout\ & ( (\Add1~113_sumout\ & \R.aluOp.ALUOpAdd~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000110000001100000011111111110000001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Add1~113_sumout\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_R.aluOp.ALUOpSub~q\,
	dataf => \ALT_INV_Add2~113_sumout\,
	combout => \Comb:vJumpAdr[28]~0_RESYN1032_BDD1033\);

-- Location: MLABCELL_X78_Y4_N6
\Comb:vJumpAdr[28]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[28]~0_combout\ = ( \R.aluCalc~q\ & ( \Add3~113_sumout\ & ( ((!\Equal4~2_combout\) # (\Selector4~1_combout\)) # (\Comb:vJumpAdr[28]~0_RESYN1032_BDD1033\) ) ) ) # ( !\R.aluCalc~q\ & ( \Add3~113_sumout\ & ( (!\Equal4~2_combout\) # 
-- (\R.aluRes\(28)) ) ) ) # ( \R.aluCalc~q\ & ( !\Add3~113_sumout\ & ( (\Equal4~2_combout\ & ((\Selector4~1_combout\) # (\Comb:vJumpAdr[28]~0_RESYN1032_BDD1033\))) ) ) ) # ( !\R.aluCalc~q\ & ( !\Add3~113_sumout\ & ( (\R.aluRes\(28) & \Equal4~2_combout\) ) ) 
-- )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000001111000000000111011111111111000011111111111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Comb:vJumpAdr[28]~0_RESYN1032_BDD1033\,
	datab => \ALT_INV_Selector4~1_combout\,
	datac => \ALT_INV_R.aluRes\(28),
	datad => \ALT_INV_Equal4~2_combout\,
	datae => \ALT_INV_R.aluCalc~q\,
	dataf => \ALT_INV_Add3~113_sumout\,
	combout => \Comb:vJumpAdr[28]~0_combout\);

-- Location: FF_X78_Y4_N7
\R.curPC[28]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[28]~0_combout\,
	asdata => \Add0~105_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(28));

-- Location: MLABCELL_X65_Y1_N48
\Mux62~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux62~14_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[8][28]~q\))) # (\R.curInst\(15) & (\RegFile[9][28]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[10][28]~q\))) # (\R.curInst\(15) & (\RegFile[11][28]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[11][28]~q\,
	datab => \ALT_INV_RegFile[9][28]~q\,
	datac => \ALT_INV_RegFile[10][28]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][28]~q\,
	combout => \Mux62~14_combout\);

-- Location: MLABCELL_X65_Y1_N36
\Mux62~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux62~1_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux62~14_combout\)))) # (\R.curInst\(17) & ((!\Mux62~14_combout\ & ((\RegFile[12][28]~q\))) # (\Mux62~14_combout\ & (\RegFile[13][28]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux62~14_combout\)))) # (\R.curInst\(17) & ((!\Mux62~14_combout\ & ((\RegFile[14][28]~q\))) # (\Mux62~14_combout\ & (\RegFile[15][28]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][28]~q\,
	datab => \ALT_INV_RegFile[15][28]~q\,
	datac => \ALT_INV_RegFile[14][28]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux62~14_combout\,
	datag => \ALT_INV_RegFile[12][28]~q\,
	combout => \Mux62~1_combout\);

-- Location: FF_X61_Y1_N44
\RegFile[6][28]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(28),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[6][28]~DUPLICATE_q\);

-- Location: LABCELL_X61_Y1_N36
\Mux62~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux62~0_combout\ = ( \RegFile[7][28]~q\ & ( \R.curInst\(15) & ( (\R.curInst\(16)) # (\RegFile[5][28]~q\) ) ) ) # ( !\RegFile[7][28]~q\ & ( \R.curInst\(15) & ( (\RegFile[5][28]~q\ & !\R.curInst\(16)) ) ) ) # ( \RegFile[7][28]~q\ & ( !\R.curInst\(15) & ( 
-- (!\R.curInst\(16) & ((\RegFile[4][28]~q\))) # (\R.curInst\(16) & (\RegFile[6][28]~DUPLICATE_q\)) ) ) ) # ( !\RegFile[7][28]~q\ & ( !\R.curInst\(15) & ( (!\R.curInst\(16) & ((\RegFile[4][28]~q\))) # (\R.curInst\(16) & (\RegFile[6][28]~DUPLICATE_q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100110011000011110011001101010101000000000101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[5][28]~q\,
	datab => \ALT_INV_RegFile[6][28]~DUPLICATE_q\,
	datac => \ALT_INV_RegFile[4][28]~q\,
	datad => \ALT_INV_R.curInst\(16),
	datae => \ALT_INV_RegFile[7][28]~q\,
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux62~0_combout\);

-- Location: LABCELL_X70_Y5_N24
\Mux62~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux62~26_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (\R.curInst\(15) & (\RegFile[1][28]~q\))) # (\R.curInst\(17) & (((\Mux62~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & ((!\R.curInst\(15) & (((\RegFile[2][28]~q\)))) # 
-- (\R.curInst\(15) & (\RegFile[3][28]~q\)))) # (\R.curInst\(17) & ((((\Mux62~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000000000111010000000000000011111111110001110111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][28]~q\,
	datab => \ALT_INV_R.curInst\(15),
	datac => \ALT_INV_RegFile[2][28]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux62~0_combout\,
	datag => \ALT_INV_RegFile[1][28]~q\,
	combout => \Mux62~26_combout\);

-- Location: LABCELL_X67_Y4_N18
\Mux62~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux62~22_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[24][28]~q\))) # (\R.curInst\(15) & (\RegFile[25][28]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & (\RegFile[26][28]~q\)) # (\R.curInst\(15) & ((\RegFile[27][28]~q\)))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001110111011101110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[25][28]~q\,
	datac => \ALT_INV_RegFile[26][28]~q\,
	datad => \ALT_INV_RegFile[27][28]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][28]~q\,
	combout => \Mux62~22_combout\);

-- Location: LABCELL_X70_Y5_N0
\Mux62~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux62~9_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux62~22_combout\)))) # (\R.curInst\(17) & ((!\Mux62~22_combout\ & ((\RegFile[28][28]~q\))) # (\Mux62~22_combout\ & (\RegFile[29][28]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux62~22_combout\)))) # (\R.curInst\(17) & ((!\Mux62~22_combout\ & ((\RegFile[30][28]~q\))) # (\Mux62~22_combout\ & (\RegFile[31][28]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][28]~q\,
	datab => \ALT_INV_RegFile[29][28]~q\,
	datac => \ALT_INV_RegFile[30][28]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux62~22_combout\,
	datag => \ALT_INV_RegFile[28][28]~q\,
	combout => \Mux62~9_combout\);

-- Location: LABCELL_X67_Y9_N48
\Mux62~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux62~18_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[16][28]~q\))) # (\R.curInst\(15) & (\RegFile[17][28]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[18][28]~q\))) # (\R.curInst\(15) & (\RegFile[19][28]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[19][28]~q\,
	datab => \ALT_INV_RegFile[17][28]~q\,
	datac => \ALT_INV_RegFile[18][28]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][28]~q\,
	combout => \Mux62~18_combout\);

-- Location: LABCELL_X70_Y5_N33
\Mux62~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux62~5_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux62~18_combout\))))) # (\R.curInst\(17) & (((!\Mux62~18_combout\ & ((\RegFile[20][28]~q\))) # (\Mux62~18_combout\ & (\RegFile[21][28]~q\))))) ) ) # ( \R.curInst\(16) & ( 
-- ((!\R.curInst\(17) & (((\Mux62~18_combout\)))) # (\R.curInst\(17) & ((!\Mux62~18_combout\ & (\RegFile[22][28]~q\)) # (\Mux62~18_combout\ & ((\RegFile[23][28]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][28]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[22][28]~q\,
	datad => \ALT_INV_RegFile[23][28]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux62~18_combout\,
	datag => \ALT_INV_RegFile[20][28]~q\,
	combout => \Mux62~5_combout\);

-- Location: LABCELL_X70_Y5_N9
\Mux62~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux62~13_combout\ = ( \Mux62~9_combout\ & ( \Mux62~5_combout\ & ( ((!\R.curInst\(18) & ((\Mux62~26_combout\))) # (\R.curInst\(18) & (\Mux62~1_combout\))) # (\R.curInst\(19)) ) ) ) # ( !\Mux62~9_combout\ & ( \Mux62~5_combout\ & ( (!\R.curInst\(18) & 
-- (((\Mux62~26_combout\) # (\R.curInst\(19))))) # (\R.curInst\(18) & (\Mux62~1_combout\ & (!\R.curInst\(19)))) ) ) ) # ( \Mux62~9_combout\ & ( !\Mux62~5_combout\ & ( (!\R.curInst\(18) & (((!\R.curInst\(19) & \Mux62~26_combout\)))) # (\R.curInst\(18) & 
-- (((\R.curInst\(19))) # (\Mux62~1_combout\))) ) ) ) # ( !\Mux62~9_combout\ & ( !\Mux62~5_combout\ & ( (!\R.curInst\(19) & ((!\R.curInst\(18) & ((\Mux62~26_combout\))) # (\R.curInst\(18) & (\Mux62~1_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000011010000000100111101001100011100110111000001111111011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux62~1_combout\,
	datab => \ALT_INV_R.curInst\(18),
	datac => \ALT_INV_R.curInst\(19),
	datad => \ALT_INV_Mux62~26_combout\,
	datae => \ALT_INV_Mux62~9_combout\,
	dataf => \ALT_INV_Mux62~5_combout\,
	combout => \Mux62~13_combout\);

-- Location: LABCELL_X73_Y5_N33
\Mux226~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux226~0_combout\ = ( \Mux62~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC\(28)))) ) ) # ( !\Mux62~13_combout\ & ( (\vAluSrc1~2_combout\ & (!\vAluSrc1~1_combout\ & \R.curPC\(28))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001000100000000000100010010001000110011001000100011001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluSrc1~2_combout\,
	datab => \ALT_INV_vAluSrc1~1_combout\,
	datad => \ALT_INV_R.curPC\(28),
	dataf => \ALT_INV_Mux62~13_combout\,
	combout => \Mux226~0_combout\);

-- Location: LABCELL_X74_Y5_N0
\ShiftRight1~27\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~27_combout\ = ( \Mux228~0_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (\Mux226~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & ((\Mux225~0_combout\))) ) ) ) # ( !\Mux228~0_combout\ & ( 
-- \NxR.aluData2[1]~17_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & (\Mux226~0_combout\)) # (\NxR.aluData2[0]~16_combout\ & ((\Mux225~0_combout\))) ) ) ) # ( \Mux228~0_combout\ & ( !\NxR.aluData2[1]~17_combout\ & ( (!\NxR.aluData2[0]~16_combout\) # 
-- (\Mux227~0_combout\) ) ) ) # ( !\Mux228~0_combout\ & ( !\NxR.aluData2[1]~17_combout\ & ( (\NxR.aluData2[0]~16_combout\ & \Mux227~0_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101101011111010111100100010011101110010001001110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datab => \ALT_INV_Mux226~0_combout\,
	datac => \ALT_INV_Mux227~0_combout\,
	datad => \ALT_INV_Mux225~0_combout\,
	datae => \ALT_INV_Mux228~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[1]~17_combout\,
	combout => \ShiftRight1~27_combout\);

-- Location: FF_X74_Y5_N1
\ShiftRight1~27_NEW_REG18\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~27_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~27_OTERM19\);

-- Location: MLABCELL_X82_Y6_N27
\ShiftRight1~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~29_combout\ = ( \R.aluData2\(3) & ( \ShiftRight1~28_OTERM23\ & ( (\ShiftRight1~27_OTERM19\) # (\R.aluData2\(2)) ) ) ) # ( !\R.aluData2\(3) & ( \ShiftRight1~28_OTERM23\ & ( (!\R.aluData2\(2) & (\ShiftRight1~25_OTERM277\)) # (\R.aluData2\(2) & 
-- ((\ShiftRight1~26_OTERM37\))) ) ) ) # ( \R.aluData2\(3) & ( !\ShiftRight1~28_OTERM23\ & ( (!\R.aluData2\(2) & \ShiftRight1~27_OTERM19\) ) ) ) # ( !\R.aluData2\(3) & ( !\ShiftRight1~28_OTERM23\ & ( (!\R.aluData2\(2) & (\ShiftRight1~25_OTERM277\)) # 
-- (\R.aluData2\(2) & ((\ShiftRight1~26_OTERM37\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101001011111001000100010001000001010010111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(2),
	datab => \ALT_INV_ShiftRight1~27_OTERM19\,
	datac => \ALT_INV_ShiftRight1~25_OTERM277\,
	datad => \ALT_INV_ShiftRight1~26_OTERM37\,
	datae => \ALT_INV_R.aluData2\(3),
	dataf => \ALT_INV_ShiftRight1~28_OTERM23\,
	combout => \ShiftRight1~29_combout\);

-- Location: MLABCELL_X82_Y7_N39
\Selector30~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector30~0_combout\ = ( \Add1~9_sumout\ & ( ((\Selector31~6_OTERM381\ & \ShiftRight1~29_combout\)) # (\R.aluOp.ALUOpAdd~q\) ) ) # ( !\Add1~9_sumout\ & ( (\Selector31~6_OTERM381\ & \ShiftRight1~29_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010101000000000101010100001111010111110000111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector31~6_OTERM381\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_ShiftRight1~29_combout\,
	dataf => \ALT_INV_Add1~9_sumout\,
	combout => \Selector30~0_combout\);

-- Location: LABCELL_X80_Y7_N24
\ShiftRight1~20\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~20_combout\ = ( \R.aluData2\(1) & ( \R.aluData1\(5) & ( (\R.aluData1\(4)) # (\R.aluData2\(0)) ) ) ) # ( !\R.aluData2\(1) & ( \R.aluData1\(5) & ( (!\R.aluData2\(0) & ((\R.aluData1\(2)))) # (\R.aluData2\(0) & (\R.aluData1\(3))) ) ) ) # ( 
-- \R.aluData2\(1) & ( !\R.aluData1\(5) & ( (!\R.aluData2\(0) & \R.aluData1\(4)) ) ) ) # ( !\R.aluData2\(1) & ( !\R.aluData1\(5) & ( (!\R.aluData2\(0) & ((\R.aluData1\(2)))) # (\R.aluData2\(0) & (\R.aluData1\(3))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000110111011000010100000101000010001101110110101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(0),
	datab => \ALT_INV_R.aluData1\(3),
	datac => \ALT_INV_R.aluData1\(4),
	datad => \ALT_INV_R.aluData1\(2),
	datae => \ALT_INV_R.aluData2\(1),
	dataf => \ALT_INV_R.aluData1\(5),
	combout => \ShiftRight1~20_combout\);

-- Location: LABCELL_X83_Y7_N30
\ShiftRight1~24\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~24_combout\ = ( \R.aluData2\(3) & ( \ShiftRight1~21_OTERM271\ & ( (!\R.aluData2\(2) & (\ShiftRight1~22_OTERM273\)) # (\R.aluData2\(2) & ((\ShiftRight1~23_OTERM275\))) ) ) ) # ( !\R.aluData2\(3) & ( \ShiftRight1~21_OTERM271\ & ( 
-- (\R.aluData2\(2)) # (\ShiftRight1~20_combout\) ) ) ) # ( \R.aluData2\(3) & ( !\ShiftRight1~21_OTERM271\ & ( (!\R.aluData2\(2) & (\ShiftRight1~22_OTERM273\)) # (\R.aluData2\(2) & ((\ShiftRight1~23_OTERM275\))) ) ) ) # ( !\R.aluData2\(3) & ( 
-- !\ShiftRight1~21_OTERM271\ & ( (\ShiftRight1~20_combout\ & !\R.aluData2\(2)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011000000110000010100000101111100111111001111110101000001011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~22_OTERM273\,
	datab => \ALT_INV_ShiftRight1~20_combout\,
	datac => \ALT_INV_R.aluData2\(2),
	datad => \ALT_INV_ShiftRight1~23_OTERM275\,
	datae => \ALT_INV_R.aluData2\(3),
	dataf => \ALT_INV_ShiftRight1~21_OTERM271\,
	combout => \ShiftRight1~24_combout\);

-- Location: LABCELL_X71_Y7_N18
\Selector30~1_RTM0405\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector30~1_RTM0405_combout\ = ( \NxR.aluData2[2]~19_combout\ & ( ((!\Mux252~0_combout\ & (\R.aluOp.ALUOpXor_OTERM355\)) # (\Mux252~0_combout\ & ((\R.aluOp.ALUOpAnd_OTERM357\)))) # (\R.aluOp.ALUOpOr_OTERM353\) ) ) # ( !\NxR.aluData2[2]~19_combout\ & ( 
-- (\Mux252~0_combout\ & ((\R.aluOp.ALUOpOr_OTERM353\) # (\R.aluOp.ALUOpXor_OTERM355\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000011100000111000001110000011101110011011111110111001101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpXor_OTERM355\,
	datab => \ALT_INV_R.aluOp.ALUOpOr_OTERM353\,
	datac => \ALT_INV_Mux252~0_combout\,
	datad => \ALT_INV_R.aluOp.ALUOpAnd_OTERM357\,
	dataf => \ALT_INV_NxR.aluData2[2]~19_combout\,
	combout => \Selector30~1_RTM0405_combout\);

-- Location: FF_X71_Y7_N19
\Selector30~1_NEW_REG402\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector30~1_RTM0405_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector30~1_OTERM403\);

-- Location: LABCELL_X83_Y7_N51
\Selector30~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector30~2_combout\ = ( \ShiftLeft0~2_OTERM221\ & ( !\Selector30~1_OTERM403\ & ( !\Selector32~3_OTERM379\ ) ) ) # ( !\ShiftLeft0~2_OTERM221\ & ( !\Selector30~1_OTERM403\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111101010101010101000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector32~3_OTERM379\,
	datae => \ALT_INV_ShiftLeft0~2_OTERM221\,
	dataf => \ALT_INV_Selector30~1_OTERM403\,
	combout => \Selector30~2_combout\);

-- Location: MLABCELL_X82_Y7_N12
\Selector30~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector30~3_combout\ = ( \Add2~9_sumout\ & ( (\Selector30~2_combout\ & (!\R.aluOp.ALUOpSub~q\ & ((!\ShiftRight0~3_combout\) # (!\Selector31~7_OTERM383\)))) ) ) # ( !\Add2~9_sumout\ & ( (\Selector30~2_combout\ & ((!\ShiftRight0~3_combout\) # 
-- (!\Selector31~7_OTERM383\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100100010001100110010001000110000001000000011000000100000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight0~3_combout\,
	datab => \ALT_INV_Selector30~2_combout\,
	datac => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datad => \ALT_INV_Selector31~7_OTERM383\,
	dataf => \ALT_INV_Add2~9_sumout\,
	combout => \Selector30~3_combout\);

-- Location: MLABCELL_X82_Y7_N42
\Selector30~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector30~4_combout\ = ( \Selector30~3_combout\ & ( ((\ShiftRight1~24_combout\ & \Selector31~5_OTERM599\)) # (\Selector30~0_combout\) ) ) # ( !\Selector30~3_combout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111111111111111111100110011001111110011001100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Selector30~0_combout\,
	datac => \ALT_INV_ShiftRight1~24_combout\,
	datad => \ALT_INV_Selector31~5_OTERM599\,
	dataf => \ALT_INV_Selector30~3_combout\,
	combout => \Selector30~4_combout\);

-- Location: FF_X82_Y7_N43
\R.aluRes[2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector30~4_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(2));

-- Location: MLABCELL_X82_Y7_N36
\vAluRes~2_RESYN1064\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~2_RESYN1064_BDD1065\ = ( \Selector31~6_OTERM381\ & ( ((\Selector31~5_OTERM599\ & \ShiftRight1~24_combout\)) # (\ShiftRight1~29_combout\) ) ) # ( !\Selector31~6_OTERM381\ & ( (\Selector31~5_OTERM599\ & \ShiftRight1~24_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000110000001100000011111111110000001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Selector31~5_OTERM599\,
	datac => \ALT_INV_ShiftRight1~24_combout\,
	datad => \ALT_INV_ShiftRight1~29_combout\,
	dataf => \ALT_INV_Selector31~6_OTERM381\,
	combout => \vAluRes~2_RESYN1064_BDD1065\);

-- Location: MLABCELL_X82_Y7_N24
\vAluRes~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~2_combout\ = ( \vAluRes~2_RESYN1064_BDD1065\ & ( \Selector30~3_combout\ & ( (\R.aluCalc~q\) # (\R.aluRes\(2)) ) ) ) # ( !\vAluRes~2_RESYN1064_BDD1065\ & ( \Selector30~3_combout\ & ( (!\R.aluCalc~q\ & (\R.aluRes\(2))) # (\R.aluCalc~q\ & 
-- (((\R.aluOp.ALUOpAdd~q\ & \Add1~9_sumout\)))) ) ) ) # ( \vAluRes~2_RESYN1064_BDD1065\ & ( !\Selector30~3_combout\ & ( (\R.aluCalc~q\) # (\R.aluRes\(2)) ) ) ) # ( !\vAluRes~2_RESYN1064_BDD1065\ & ( !\Selector30~3_combout\ & ( (\R.aluCalc~q\) # 
-- (\R.aluRes\(2)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010111111111010101011111111101010101000000110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluRes\(2),
	datab => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datac => \ALT_INV_Add1~9_sumout\,
	datad => \ALT_INV_R.aluCalc~q\,
	datae => \ALT_INV_vAluRes~2_RESYN1064_BDD1065\,
	dataf => \ALT_INV_Selector30~3_combout\,
	combout => \vAluRes~2_combout\);

-- Location: MLABCELL_X78_Y7_N0
\Comb:vJumpAdr[2]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[2]~0_combout\ = ( \Add3~9_sumout\ & ( (!\Equal4~2_combout\) # (\vAluRes~2_combout\) ) ) # ( !\Add3~9_sumout\ & ( (\Equal4~2_combout\ & \vAluRes~2_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101000001010000010110101111101011111010111110101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Equal4~2_combout\,
	datac => \ALT_INV_vAluRes~2_combout\,
	dataf => \ALT_INV_Add3~9_sumout\,
	combout => \Comb:vJumpAdr[2]~0_combout\);

-- Location: FF_X78_Y7_N1
\R.curPC[2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[2]~0_combout\,
	asdata => \Add0~1_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(2));

-- Location: MLABCELL_X82_Y7_N15
\R.regWriteData[2]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.regWriteData[2]~feeder_combout\ = ( \Add0~1_sumout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_Add0~1_sumout\,
	combout => \R.regWriteData[2]~feeder_combout\);

-- Location: IOIBUF_X89_Y13_N21
\avm_d_readdata[26]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(26),
	o => \avm_d_readdata[26]~input_o\);

-- Location: LABCELL_X83_Y5_N6
\Comb:vRegWriteData[2]~0_RESYN1082\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[2]~0_RESYN1082_BDD1083\ = ( \Mux222~0_combout\ & ( \R.memToReg~q\ & ( \avm_d_readdata[26]~input_o\ ) ) ) # ( \Mux222~0_combout\ & ( !\R.memToReg~q\ & ( (!\R.aluCalc~q\ & ((\R.aluRes\(2)))) # (\R.aluCalc~q\ & (\Selector31~5_OTERM599\)) 
-- ) ) ) # ( !\Mux222~0_combout\ & ( !\R.memToReg~q\ & ( (!\R.aluCalc~q\ & ((\R.aluRes\(2)))) # (\R.aluCalc~q\ & (\Selector31~5_OTERM599\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001101100011011000110110001101100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluCalc~q\,
	datab => \ALT_INV_Selector31~5_OTERM599\,
	datac => \ALT_INV_R.aluRes\(2),
	datad => \ALT_INV_avm_d_readdata[26]~input_o\,
	datae => \ALT_INV_Mux222~0_combout\,
	dataf => \ALT_INV_R.memToReg~q\,
	combout => \Comb:vRegWriteData[2]~0_RESYN1082_BDD1083\);

-- Location: MLABCELL_X82_Y7_N54
\Comb:vRegWriteData[2]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[2]~0_combout\ = ( \R.aluCalc~q\ & ( \Comb:vRegWriteData[2]~0_RESYN1082_BDD1083\ & ( ((!\Selector30~3_combout\) # ((\Selector30~0_combout\) # (\R.memToReg~q\))) # (\ShiftRight1~24_combout\) ) ) ) # ( !\R.aluCalc~q\ & ( 
-- \Comb:vRegWriteData[2]~0_RESYN1082_BDD1083\ ) ) # ( \R.aluCalc~q\ & ( !\Comb:vRegWriteData[2]~0_RESYN1082_BDD1083\ & ( (!\R.memToReg~q\ & ((!\Selector30~3_combout\) # (\Selector30~0_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110000001111000011111111111111111101111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~24_combout\,
	datab => \ALT_INV_Selector30~3_combout\,
	datac => \ALT_INV_R.memToReg~q\,
	datad => \ALT_INV_Selector30~0_combout\,
	datae => \ALT_INV_R.aluCalc~q\,
	dataf => \ALT_INV_Comb:vRegWriteData[2]~0_RESYN1082_BDD1083\,
	combout => \Comb:vRegWriteData[2]~0_combout\);

-- Location: FF_X82_Y7_N17
\R.regWriteData[2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \R.regWriteData[2]~feeder_combout\,
	asdata => \Comb:vRegWriteData[2]~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(2));

-- Location: FF_X66_Y9_N2
\RegFile[2][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(2),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~4_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[2][2]~q\);

-- Location: LABCELL_X70_Y9_N33
\Mux120~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux120~0_combout\ = ( \R.curInst\(20) & ( \R.curInst\(21) & ( \RegFile[7][2]~q\ ) ) ) # ( !\R.curInst\(20) & ( \R.curInst\(21) & ( \RegFile[6][2]~q\ ) ) ) # ( \R.curInst\(20) & ( !\R.curInst\(21) & ( \RegFile[5][2]~q\ ) ) ) # ( !\R.curInst\(20) & ( 
-- !\R.curInst\(21) & ( \RegFile[4][2]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111001100110011001101010101010101010000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[6][2]~q\,
	datab => \ALT_INV_RegFile[5][2]~q\,
	datac => \ALT_INV_RegFile[7][2]~q\,
	datad => \ALT_INV_RegFile[4][2]~q\,
	datae => \ALT_INV_R.curInst\(20),
	dataf => \ALT_INV_R.curInst\(21),
	combout => \Mux120~0_combout\);

-- Location: LABCELL_X71_Y7_N6
\Mux120~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux120~26_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (\R.curInst\(20) & (\RegFile[1][2]~q\))) # (\R.curInst\(22) & ((((\Mux120~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (\RegFile[2][2]~q\)) # 
-- (\R.curInst\(20) & (((\RegFile[3][2]~q\)))))) # (\R.curInst\(22) & ((((\Mux120~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010000000100000010000100110000110111001101110011101101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(20),
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[2][2]~q\,
	datad => \ALT_INV_RegFile[3][2]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux120~0_combout\,
	datag => \ALT_INV_RegFile[1][2]~q\,
	combout => \Mux120~26_combout\);

-- Location: FF_X66_Y10_N8
\RegFile[14][2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(2),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~10_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[14][2]~q\);

-- Location: LABCELL_X66_Y7_N12
\Mux120~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux120~14_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[8][2]~q\))) # (\R.curInst\(20) & (\RegFile[9][2]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[10][2]~q\))) # (\R.curInst\(20) & (\RegFile[11][2]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][2]~q\,
	datab => \ALT_INV_RegFile[11][2]~q\,
	datac => \ALT_INV_RegFile[10][2]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][2]~q\,
	combout => \Mux120~14_combout\);

-- Location: LABCELL_X71_Y7_N36
\Mux120~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux120~1_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux120~14_combout\)))) # (\R.curInst\(22) & ((!\Mux120~14_combout\ & ((\RegFile[12][2]~q\))) # (\Mux120~14_combout\ & (\RegFile[13][2]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux120~14_combout\)))) # (\R.curInst\(22) & ((!\Mux120~14_combout\ & ((\RegFile[14][2]~q\))) # (\Mux120~14_combout\ & (\RegFile[15][2]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][2]~q\,
	datab => \ALT_INV_RegFile[15][2]~q\,
	datac => \ALT_INV_RegFile[14][2]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux120~14_combout\,
	datag => \ALT_INV_RegFile[12][2]~q\,
	combout => \Mux120~1_combout\);

-- Location: LABCELL_X68_Y8_N9
\Mux120~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux120~18_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[16][2]~q\))) # (\R.curInst\(20) & (\RegFile[17][2]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & (\RegFile[18][2]~q\)) # (\R.curInst\(20) & ((\RegFile[19][2]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[17][2]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[18][2]~q\,
	datad => \ALT_INV_RegFile[19][2]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][2]~q\,
	combout => \Mux120~18_combout\);

-- Location: MLABCELL_X72_Y8_N0
\Mux120~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux120~5_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux120~18_combout\)))) # (\R.curInst\(22) & ((!\Mux120~18_combout\ & ((\RegFile[20][2]~q\))) # (\Mux120~18_combout\ & (\RegFile[21][2]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux120~18_combout\)))) # (\R.curInst\(22) & ((!\Mux120~18_combout\ & ((\RegFile[22][2]~q\))) # (\Mux120~18_combout\ & (\RegFile[23][2]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][2]~q\,
	datab => \ALT_INV_RegFile[23][2]~q\,
	datac => \ALT_INV_RegFile[22][2]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux120~18_combout\,
	datag => \ALT_INV_RegFile[20][2]~q\,
	combout => \Mux120~5_combout\);

-- Location: LABCELL_X70_Y10_N42
\Mux120~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux120~22_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[24][2]~q\))) # (\R.curInst\(20) & (\RegFile[25][2]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & (\RegFile[26][2]~q\)) # (\R.curInst\(20) & ((\RegFile[27][2]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[25][2]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[26][2]~q\,
	datad => \ALT_INV_RegFile[27][2]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][2]~q\,
	combout => \Mux120~22_combout\);

-- Location: LABCELL_X70_Y10_N51
\Mux120~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux120~9_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux120~22_combout\))))) # (\R.curInst\(22) & (((!\Mux120~22_combout\ & ((\RegFile[28][2]~q\))) # (\Mux120~22_combout\ & (\RegFile[29][2]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux120~22_combout\)))) # (\R.curInst\(22) & ((!\Mux120~22_combout\ & (\RegFile[30][2]~q\)) # (\Mux120~22_combout\ & ((\RegFile[31][2]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[29][2]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[30][2]~q\,
	datad => \ALT_INV_RegFile[31][2]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux120~22_combout\,
	datag => \ALT_INV_RegFile[28][2]~q\,
	combout => \Mux120~9_combout\);

-- Location: LABCELL_X71_Y7_N48
\Mux120~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux120~13_combout\ = ( \Mux120~5_combout\ & ( \Mux120~9_combout\ & ( ((!\R.curInst\(23) & (\Mux120~26_combout\)) # (\R.curInst\(23) & ((\Mux120~1_combout\)))) # (\R.curInst\(24)) ) ) ) # ( !\Mux120~5_combout\ & ( \Mux120~9_combout\ & ( (!\R.curInst\(24) 
-- & ((!\R.curInst\(23) & (\Mux120~26_combout\)) # (\R.curInst\(23) & ((\Mux120~1_combout\))))) # (\R.curInst\(24) & (\R.curInst\(23))) ) ) ) # ( \Mux120~5_combout\ & ( !\Mux120~9_combout\ & ( (!\R.curInst\(24) & ((!\R.curInst\(23) & (\Mux120~26_combout\)) # 
-- (\R.curInst\(23) & ((\Mux120~1_combout\))))) # (\R.curInst\(24) & (!\R.curInst\(23))) ) ) ) # ( !\Mux120~5_combout\ & ( !\Mux120~9_combout\ & ( (!\R.curInst\(24) & ((!\R.curInst\(23) & (\Mux120~26_combout\)) # (\R.curInst\(23) & ((\Mux120~1_combout\))))) 
-- ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000100000101010010011000110111000011001001110110101110101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(24),
	datab => \ALT_INV_R.curInst\(23),
	datac => \ALT_INV_Mux120~26_combout\,
	datad => \ALT_INV_Mux120~1_combout\,
	datae => \ALT_INV_Mux120~5_combout\,
	dataf => \ALT_INV_Mux120~9_combout\,
	combout => \Mux120~13_combout\);

-- Location: LABCELL_X71_Y7_N27
\NxR.aluData2[2]~19\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[2]~19_combout\ = ( \Mux120~13_combout\ & ( (!\vAluSrc2~1_combout\) # ((\Equal4~1_combout\ & \Mux152~0_combout\)) ) ) # ( !\Mux120~13_combout\ & ( (\Equal4~1_combout\ & (\Mux152~0_combout\ & \vAluSrc2~1_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000101000000000000010111111111000001011111111100000101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Equal4~1_combout\,
	datac => \ALT_INV_Mux152~0_combout\,
	datad => \ALT_INV_vAluSrc2~1_combout\,
	dataf => \ALT_INV_Mux120~13_combout\,
	combout => \NxR.aluData2[2]~19_combout\);

-- Location: LABCELL_X71_Y7_N57
\Selector32~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector32~3_combout\ = ( \R.aluOp.ALUOpSLL_OTERM359\ & ( (!\NxR.aluData2[2]~19_combout\ & (!\NxR.aluData2[4]~20_combout\ & !\NxR.aluData2[3]~18_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000010100000000000001010000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_NxR.aluData2[2]~19_combout\,
	datac => \ALT_INV_NxR.aluData2[4]~20_combout\,
	datad => \ALT_INV_NxR.aluData2[3]~18_combout\,
	dataf => \ALT_INV_R.aluOp.ALUOpSLL_OTERM359\,
	combout => \Selector32~3_combout\);

-- Location: FF_X71_Y7_N58
\Selector32~3_NEW_REG378\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector32~3_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector32~3_OTERM379\);

-- Location: MLABCELL_X72_Y7_N30
\Selector31~2_RTM0401\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector31~2_RTM0401_combout\ = ( \R.aluOp.ALUOpAnd_OTERM357\ & ( (!\Mux253~0_combout\ & (\NxR.aluData2[1]~17_combout\ & ((\R.aluOp.ALUOpXor_OTERM355\) # (\R.aluOp.ALUOpOr_OTERM353\)))) # (\Mux253~0_combout\ & (((\R.aluOp.ALUOpXor_OTERM355\) # 
-- (\R.aluOp.ALUOpOr_OTERM353\)) # (\NxR.aluData2[1]~17_combout\))) ) ) # ( !\R.aluOp.ALUOpAnd_OTERM357\ & ( (!\R.aluOp.ALUOpOr_OTERM353\ & (\R.aluOp.ALUOpXor_OTERM355\ & (!\Mux253~0_combout\ $ (!\NxR.aluData2[1]~17_combout\)))) # (\R.aluOp.ALUOpOr_OTERM353\ 
-- & (((\NxR.aluData2[1]~17_combout\)) # (\Mux253~0_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000011101100111000001110110011100010111011101110001011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux253~0_combout\,
	datab => \ALT_INV_NxR.aluData2[1]~17_combout\,
	datac => \ALT_INV_R.aluOp.ALUOpOr_OTERM353\,
	datad => \ALT_INV_R.aluOp.ALUOpXor_OTERM355\,
	dataf => \ALT_INV_R.aluOp.ALUOpAnd_OTERM357\,
	combout => \Selector31~2_RTM0401_combout\);

-- Location: FF_X72_Y7_N31
\Selector31~2_NEW_REG398\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector31~2_RTM0401_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector31~2_OTERM399\);

-- Location: LABCELL_X83_Y7_N36
\Selector31~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector31~3_combout\ = ( !\Selector31~2_OTERM399\ & ( \ShiftLeft0~1_OTERM255\ & ( !\Selector32~3_OTERM379\ ) ) ) # ( !\Selector31~2_OTERM399\ & ( !\ShiftLeft0~1_OTERM255\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111000000000000000011110000111100000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Selector32~3_OTERM379\,
	datae => \ALT_INV_Selector31~2_OTERM399\,
	dataf => \ALT_INV_ShiftLeft0~1_OTERM255\,
	combout => \Selector31~3_combout\);

-- Location: LABCELL_X81_Y9_N27
\Selector31~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector31~4_combout\ = ( \Add2~5_sumout\ & ( \Add1~5_sumout\ & ( (\Selector31~3_combout\ & (!\R.aluOp.ALUOpAdd~q\ & !\R.aluOp.ALUOpSub~q\)) ) ) ) # ( !\Add2~5_sumout\ & ( \Add1~5_sumout\ & ( (\Selector31~3_combout\ & !\R.aluOp.ALUOpAdd~q\) ) ) ) # ( 
-- \Add2~5_sumout\ & ( !\Add1~5_sumout\ & ( (\Selector31~3_combout\ & !\R.aluOp.ALUOpSub~q\) ) ) ) # ( !\Add2~5_sumout\ & ( !\Add1~5_sumout\ & ( \Selector31~3_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101010101010000000001010000010100000101000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector31~3_combout\,
	datac => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datad => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datae => \ALT_INV_Add2~5_sumout\,
	dataf => \ALT_INV_Add1~5_sumout\,
	combout => \Selector31~4_combout\);

-- Location: LABCELL_X83_Y5_N42
\Comb:vJumpAdr[1]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[1]~0_combout\ = ( \R.aluCalc~q\ & ( \Add3~5_sumout\ & ( (!\Selector31~4_combout\) # ((!\Equal4~2_combout\) # (\Selector31~1_combout\)) ) ) ) # ( !\R.aluCalc~q\ & ( \Add3~5_sumout\ & ( (!\Equal4~2_combout\) # (\R.aluRes\(1)) ) ) ) # ( 
-- \R.aluCalc~q\ & ( !\Add3~5_sumout\ & ( (\Equal4~2_combout\ & ((!\Selector31~4_combout\) # (\Selector31~1_combout\))) ) ) ) # ( !\R.aluCalc~q\ & ( !\Add3~5_sumout\ & ( (\R.aluRes\(1) & \Equal4~2_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110011000000001010111111111111001100111111111110101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector31~4_combout\,
	datab => \ALT_INV_R.aluRes\(1),
	datac => \ALT_INV_Selector31~1_combout\,
	datad => \ALT_INV_Equal4~2_combout\,
	datae => \ALT_INV_R.aluCalc~q\,
	dataf => \ALT_INV_Add3~5_sumout\,
	combout => \Comb:vJumpAdr[1]~0_combout\);

-- Location: FF_X83_Y5_N43
\R.curPC[1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[1]~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(1));

-- Location: LABCELL_X70_Y9_N24
\Mux89~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux89~0_combout\ = ( \R.curInst\(16) & ( \R.curInst\(15) & ( \RegFile[7][1]~q\ ) ) ) # ( !\R.curInst\(16) & ( \R.curInst\(15) & ( \RegFile[5][1]~q\ ) ) ) # ( \R.curInst\(16) & ( !\R.curInst\(15) & ( \RegFile[6][1]~q\ ) ) ) # ( !\R.curInst\(16) & ( 
-- !\R.curInst\(15) & ( \RegFile[4][1]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110011000011110000111101010101010101010000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[5][1]~q\,
	datab => \ALT_INV_RegFile[4][1]~q\,
	datac => \ALT_INV_RegFile[6][1]~q\,
	datad => \ALT_INV_RegFile[7][1]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	combout => \Mux89~0_combout\);

-- Location: LABCELL_X70_Y9_N48
\Mux89~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux89~26_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((\RegFile[1][1]~q\ & (\R.curInst\(15)))))) # (\R.curInst\(17) & ((((\Mux89~0_combout\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & ((!\R.curInst\(15) & (((\RegFile[2][1]~q\)))) # 
-- (\R.curInst\(15) & (\RegFile[3][1]~q\)))) # (\R.curInst\(17) & ((((\Mux89~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001010000010100010001001010101010111110101111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[3][1]~q\,
	datac => \ALT_INV_RegFile[2][1]~q\,
	datad => \ALT_INV_R.curInst\(15),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux89~0_combout\,
	datag => \ALT_INV_RegFile[1][1]~q\,
	combout => \Mux89~26_combout\);

-- Location: LABCELL_X70_Y8_N24
\Mux89~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux89~22_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & ((\RegFile[24][1]~q\))) # (\R.curInst\(15) & (\RegFile[25][1]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & ((\RegFile[26][1]~q\))) # (\R.curInst\(15) & (\RegFile[27][1]~q\)))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[27][1]~q\,
	datab => \ALT_INV_RegFile[25][1]~q\,
	datac => \ALT_INV_RegFile[26][1]~q\,
	datad => \ALT_INV_R.curInst\(17),
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[24][1]~q\,
	combout => \Mux89~22_combout\);

-- Location: LABCELL_X70_Y8_N15
\Mux89~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux89~9_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & (((\Mux89~22_combout\)))) # (\R.curInst\(17) & ((!\Mux89~22_combout\ & (\RegFile[28][1]~q\)) # (\Mux89~22_combout\ & ((\RegFile[29][1]~q\)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- ((((\Mux89~22_combout\))))) # (\R.curInst\(17) & (((!\Mux89~22_combout\ & ((\RegFile[30][1]~q\))) # (\Mux89~22_combout\ & (\RegFile[31][1]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111001100111111111101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][1]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[30][1]~q\,
	datad => \ALT_INV_RegFile[29][1]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux89~22_combout\,
	datag => \ALT_INV_RegFile[28][1]~q\,
	combout => \Mux89~9_combout\);

-- Location: LABCELL_X63_Y8_N24
\Mux89~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux89~14_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & (((!\R.curInst\(15) & ((\RegFile[8][1]~q\))) # (\R.curInst\(15) & (\RegFile[9][1]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( ((!\R.curInst\(17) & 
-- ((!\R.curInst\(15) & (\RegFile[10][1]~q\)) # (\R.curInst\(15) & ((\RegFile[11][1]~q\))))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][1]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[10][1]~q\,
	datad => \ALT_INV_RegFile[11][1]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[8][1]~q\,
	combout => \Mux89~14_combout\);

-- Location: FF_X66_Y7_N35
\RegFile[12][1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[12][1]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][1]~q\);

-- Location: LABCELL_X63_Y8_N39
\Mux89~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux89~1_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux89~14_combout\))))) # (\R.curInst\(17) & (((!\Mux89~14_combout\ & ((\RegFile[12][1]~q\))) # (\Mux89~14_combout\ & (\RegFile[13][1]~q\))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) 
-- & ((((\Mux89~14_combout\))))) # (\R.curInst\(17) & (((!\Mux89~14_combout\ & (\RegFile[14][1]~q\)) # (\Mux89~14_combout\ & ((\RegFile[15][1]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110111011101110111010101011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[13][1]~q\,
	datac => \ALT_INV_RegFile[14][1]~q\,
	datad => \ALT_INV_RegFile[15][1]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux89~14_combout\,
	datag => \ALT_INV_RegFile[12][1]~q\,
	combout => \Mux89~1_combout\);

-- Location: LABCELL_X70_Y4_N18
\Mux89~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux89~18_combout\ = ( !\R.curInst\(16) & ( ((!\R.curInst\(17) & ((!\R.curInst\(15) & (\RegFile[16][1]~q\)) # (\R.curInst\(15) & ((\RegFile[17][1]~q\))))) # (\R.curInst\(17) & (((\R.curInst\(15)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) & 
-- (((!\R.curInst\(15) & ((\RegFile[18][1]~q\))) # (\R.curInst\(15) & (\RegFile[19][1]~q\))))) # (\R.curInst\(17) & ((((\R.curInst\(15)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110000110011111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[19][1]~q\,
	datab => \ALT_INV_R.curInst\(17),
	datac => \ALT_INV_RegFile[18][1]~q\,
	datad => \ALT_INV_RegFile[17][1]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_R.curInst\(15),
	datag => \ALT_INV_RegFile[16][1]~q\,
	combout => \Mux89~18_combout\);

-- Location: LABCELL_X70_Y4_N42
\Mux89~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux89~5_combout\ = ( !\R.curInst\(16) & ( (!\R.curInst\(17) & ((((\Mux89~18_combout\))))) # (\R.curInst\(17) & (((!\Mux89~18_combout\ & (\RegFile[20][1]~q\)) # (\Mux89~18_combout\ & ((\RegFile[21][1]~q\)))))) ) ) # ( \R.curInst\(16) & ( (!\R.curInst\(17) 
-- & ((((\Mux89~18_combout\))))) # (\R.curInst\(17) & (((!\Mux89~18_combout\ & ((\RegFile[22][1]~q\))) # (\Mux89~18_combout\ & (\RegFile[23][1]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110101010111111111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(17),
	datab => \ALT_INV_RegFile[23][1]~q\,
	datac => \ALT_INV_RegFile[22][1]~q\,
	datad => \ALT_INV_RegFile[21][1]~q\,
	datae => \ALT_INV_R.curInst\(16),
	dataf => \ALT_INV_Mux89~18_combout\,
	datag => \ALT_INV_RegFile[20][1]~q\,
	combout => \Mux89~5_combout\);

-- Location: LABCELL_X71_Y8_N48
\Mux89~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux89~13_combout\ = ( \Mux89~1_combout\ & ( \Mux89~5_combout\ & ( (!\R.curInst\(18) & (((\Mux89~26_combout\)) # (\R.curInst\(19)))) # (\R.curInst\(18) & ((!\R.curInst\(19)) # ((\Mux89~9_combout\)))) ) ) ) # ( !\Mux89~1_combout\ & ( \Mux89~5_combout\ & ( 
-- (!\R.curInst\(18) & (((\Mux89~26_combout\)) # (\R.curInst\(19)))) # (\R.curInst\(18) & (\R.curInst\(19) & ((\Mux89~9_combout\)))) ) ) ) # ( \Mux89~1_combout\ & ( !\Mux89~5_combout\ & ( (!\R.curInst\(18) & (!\R.curInst\(19) & (\Mux89~26_combout\))) # 
-- (\R.curInst\(18) & ((!\R.curInst\(19)) # ((\Mux89~9_combout\)))) ) ) ) # ( !\Mux89~1_combout\ & ( !\Mux89~5_combout\ & ( (!\R.curInst\(18) & (!\R.curInst\(19) & (\Mux89~26_combout\))) # (\R.curInst\(18) & (\R.curInst\(19) & ((\Mux89~9_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000100000011001010011000101110100101010001110110110111001111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(18),
	datab => \ALT_INV_R.curInst\(19),
	datac => \ALT_INV_Mux89~26_combout\,
	datad => \ALT_INV_Mux89~9_combout\,
	datae => \ALT_INV_Mux89~1_combout\,
	dataf => \ALT_INV_Mux89~5_combout\,
	combout => \Mux89~13_combout\);

-- Location: MLABCELL_X72_Y7_N18
\Mux253~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux253~0_combout\ = ( \Mux89~13_combout\ & ( (!\vAluSrc1~1_combout\ & ((!\vAluSrc1~2_combout\) # (\R.curPC\(1)))) ) ) # ( !\Mux89~13_combout\ & ( (!\vAluSrc1~1_combout\ & (\R.curPC\(1) & \vAluSrc1~2_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000001100000000000000110011001100000011001100110000001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_vAluSrc1~1_combout\,
	datac => \ALT_INV_R.curPC\(1),
	datad => \ALT_INV_vAluSrc1~2_combout\,
	dataf => \ALT_INV_Mux89~13_combout\,
	combout => \Mux253~0_combout\);

-- Location: MLABCELL_X72_Y7_N42
\ShiftLeft0~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~5_combout\ = ( \NxR.aluData2[0]~16_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( \Mux253~0_combout\ ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( \Mux252~0_combout\ ) ) ) # ( \NxR.aluData2[0]~16_combout\ & ( 
-- !\NxR.aluData2[1]~17_combout\ & ( \Mux251~0_combout\ ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( !\NxR.aluData2[1]~17_combout\ & ( \Mux250~0_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000000001111111100110011001100110101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux253~0_combout\,
	datab => \ALT_INV_Mux252~0_combout\,
	datac => \ALT_INV_Mux250~0_combout\,
	datad => \ALT_INV_Mux251~0_combout\,
	datae => \ALT_INV_NxR.aluData2[0]~16_combout\,
	dataf => \ALT_INV_NxR.aluData2[1]~17_combout\,
	combout => \ShiftLeft0~5_combout\);

-- Location: FF_X72_Y7_N43
\ShiftLeft0~5_NEW_REG202\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftLeft0~5_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftLeft0~5_OTERM203\);

-- Location: MLABCELL_X72_Y5_N12
\Selector28~1_RTM0389\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector28~1_RTM0389_combout\ = ( \Mux250~0_combout\ & ( ((!\NxR.aluData2[4]~20_combout\ & (\R.aluOp.ALUOpXor_OTERM355\)) # (\NxR.aluData2[4]~20_combout\ & ((\R.aluOp.ALUOpAnd_OTERM357\)))) # (\R.aluOp.ALUOpOr_OTERM353\) ) ) # ( !\Mux250~0_combout\ & ( 
-- (\NxR.aluData2[4]~20_combout\ & ((\R.aluOp.ALUOpXor_OTERM355\) # (\R.aluOp.ALUOpOr_OTERM353\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000011100000111000001110000011101110101011111110111010101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpOr_OTERM353\,
	datab => \ALT_INV_R.aluOp.ALUOpXor_OTERM355\,
	datac => \ALT_INV_NxR.aluData2[4]~20_combout\,
	datad => \ALT_INV_R.aluOp.ALUOpAnd_OTERM357\,
	dataf => \ALT_INV_Mux250~0_combout\,
	combout => \Selector28~1_RTM0389_combout\);

-- Location: FF_X72_Y5_N13
\Selector28~1_NEW_REG386\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector28~1_RTM0389_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector28~1_OTERM387\);

-- Location: LABCELL_X75_Y8_N30
\Selector28~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector28~2_combout\ = ( !\Selector28~1_OTERM387\ & ( (!\Selector27~0_OTERM385\) # ((!\ShiftLeft0~4_OTERM237\ & ((!\ShiftLeft0~5_OTERM203\) # (\ShiftRight0~7_OTERM233DUPLICATE_q\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1110110011111100111011001111110000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~5_OTERM203\,
	datab => \ALT_INV_Selector27~0_OTERM385\,
	datac => \ALT_INV_ShiftLeft0~4_OTERM237\,
	datad => \ALT_INV_ShiftRight0~7_OTERM233DUPLICATE_q\,
	dataf => \ALT_INV_Selector28~1_OTERM387\,
	combout => \Selector28~2_combout\);

-- Location: LABCELL_X73_Y7_N0
\ShiftRight1~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~6_combout\ = ( \Mux247~0_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( (\NxR.aluData2[0]~16_combout\) # (\Mux248~0_combout\) ) ) ) # ( !\Mux247~0_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( (\Mux248~0_combout\ & 
-- !\NxR.aluData2[0]~16_combout\) ) ) ) # ( \Mux247~0_combout\ & ( !\NxR.aluData2[1]~17_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & ((\Mux250~0_combout\))) # (\NxR.aluData2[0]~16_combout\ & (\Mux249~0_combout\)) ) ) ) # ( !\Mux247~0_combout\ & ( 
-- !\NxR.aluData2[1]~17_combout\ & ( (!\NxR.aluData2[0]~16_combout\ & ((\Mux250~0_combout\))) # (\NxR.aluData2[0]~16_combout\ & (\Mux249~0_combout\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001101010101001100110101010100001111000000000000111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux249~0_combout\,
	datab => \ALT_INV_Mux250~0_combout\,
	datac => \ALT_INV_Mux248~0_combout\,
	datad => \ALT_INV_NxR.aluData2[0]~16_combout\,
	datae => \ALT_INV_Mux247~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[1]~17_combout\,
	combout => \ShiftRight1~6_combout\);

-- Location: FF_X73_Y7_N1
\ShiftRight1~6_NEW_REG196\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~6_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~6_OTERM197\);

-- Location: LABCELL_X74_Y8_N12
\ShiftRight1~40\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~40_combout\ = ( \ShiftRight1~7_OTERM259\ & ( \ShiftRight1~0_OTERM257\ & ( ((!\R.aluData2\(3) & (\ShiftRight1~6_OTERM197\)) # (\R.aluData2\(3) & ((\ShiftRight1~8_OTERM261\)))) # (\R.aluData2\(2)) ) ) ) # ( !\ShiftRight1~7_OTERM259\ & ( 
-- \ShiftRight1~0_OTERM257\ & ( (!\R.aluData2\(2) & ((!\R.aluData2\(3) & (\ShiftRight1~6_OTERM197\)) # (\R.aluData2\(3) & ((\ShiftRight1~8_OTERM261\))))) # (\R.aluData2\(2) & (\R.aluData2\(3))) ) ) ) # ( \ShiftRight1~7_OTERM259\ & ( !\ShiftRight1~0_OTERM257\ 
-- & ( (!\R.aluData2\(2) & ((!\R.aluData2\(3) & (\ShiftRight1~6_OTERM197\)) # (\R.aluData2\(3) & ((\ShiftRight1~8_OTERM261\))))) # (\R.aluData2\(2) & (!\R.aluData2\(3))) ) ) ) # ( !\ShiftRight1~7_OTERM259\ & ( !\ShiftRight1~0_OTERM257\ & ( (!\R.aluData2\(2) 
-- & ((!\R.aluData2\(3) & (\ShiftRight1~6_OTERM197\)) # (\R.aluData2\(3) & ((\ShiftRight1~8_OTERM261\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000100000101010010011000110111000011001001110110101110101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(2),
	datab => \ALT_INV_R.aluData2\(3),
	datac => \ALT_INV_ShiftRight1~6_OTERM197\,
	datad => \ALT_INV_ShiftRight1~8_OTERM261\,
	datae => \ALT_INV_ShiftRight1~7_OTERM259\,
	dataf => \ALT_INV_ShiftRight1~0_OTERM257\,
	combout => \ShiftRight1~40_combout\);

-- Location: LABCELL_X74_Y8_N18
\ShiftRight0~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight0~6_combout\ = ( \ShiftRight1~2_OTERM49\ & ( (!\R.aluData2\(2) & ((!\R.aluData2\(3) & ((\ShiftRight1~1_OTERM33\))) # (\R.aluData2\(3) & (\ShiftRight1~3_OTERM13\)))) # (\R.aluData2\(2) & (!\R.aluData2\(3))) ) ) # ( !\ShiftRight1~2_OTERM49\ & ( 
-- (!\R.aluData2\(2) & ((!\R.aluData2\(3) & ((\ShiftRight1~1_OTERM33\))) # (\R.aluData2\(3) & (\ShiftRight1~3_OTERM13\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001010001010000000101000101001000110110011100100011011001110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(2),
	datab => \ALT_INV_R.aluData2\(3),
	datac => \ALT_INV_ShiftRight1~3_OTERM13\,
	datad => \ALT_INV_ShiftRight1~1_OTERM33\,
	dataf => \ALT_INV_ShiftRight1~2_OTERM49\,
	combout => \ShiftRight0~6_combout\);

-- Location: LABCELL_X75_Y8_N0
\Selector28~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector28~3_combout\ = ( \ShiftRight1~40_combout\ & ( \ShiftRight0~6_combout\ & ( (!\Selector31~7_OTERM383\ & (!\Selector31~5_OTERM599\ & \Selector28~2_combout\)) ) ) ) # ( !\ShiftRight1~40_combout\ & ( \ShiftRight0~6_combout\ & ( 
-- (!\Selector31~7_OTERM383\ & \Selector28~2_combout\) ) ) ) # ( \ShiftRight1~40_combout\ & ( !\ShiftRight0~6_combout\ & ( (!\Selector31~5_OTERM599\ & \Selector28~2_combout\) ) ) ) # ( !\ShiftRight1~40_combout\ & ( !\ShiftRight0~6_combout\ & ( 
-- \Selector28~2_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111000000001111000000000000110011000000000011000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Selector31~7_OTERM383\,
	datac => \ALT_INV_Selector31~5_OTERM599\,
	datad => \ALT_INV_Selector28~2_combout\,
	datae => \ALT_INV_ShiftRight1~40_combout\,
	dataf => \ALT_INV_ShiftRight0~6_combout\,
	combout => \Selector28~3_combout\);

-- Location: LABCELL_X80_Y8_N39
\Selector28~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector28~0_combout\ = ( \Add2~17_sumout\ & ( \Add1~17_sumout\ & ( (\R.aluOp.ALUOpSub~q\) # (\R.aluOp.ALUOpAdd~q\) ) ) ) # ( !\Add2~17_sumout\ & ( \Add1~17_sumout\ & ( \R.aluOp.ALUOpAdd~q\ ) ) ) # ( \Add2~17_sumout\ & ( !\Add1~17_sumout\ & ( 
-- \R.aluOp.ALUOpSub~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000111100110011001100110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datac => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datae => \ALT_INV_Add2~17_sumout\,
	dataf => \ALT_INV_Add1~17_sumout\,
	combout => \Selector28~0_combout\);

-- Location: LABCELL_X80_Y6_N15
\Selector28~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector28~4_combout\ = ( \Selector28~0_combout\ ) # ( !\Selector28~0_combout\ & ( (!\Selector28~3_combout\) # ((\Selector31~6_OTERM381\ & \ShiftRight1~39_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111100000011111111110000001111111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Selector31~6_OTERM381\,
	datac => \ALT_INV_ShiftRight1~39_combout\,
	datad => \ALT_INV_Selector28~3_combout\,
	dataf => \ALT_INV_Selector28~0_combout\,
	combout => \Selector28~4_combout\);

-- Location: FF_X80_Y6_N16
\R.aluRes[4]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector28~4_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes[4]~DUPLICATE_q\);

-- Location: LABCELL_X80_Y8_N21
\vAluRes~4_RESYN1068\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~4_RESYN1068_BDD1069\ = ( \ShiftRight1~39_combout\ & ( ((\Add2~17_sumout\ & \R.aluOp.ALUOpSub~q\)) # (\Selector31~6_OTERM381\) ) ) # ( !\ShiftRight1~39_combout\ & ( (\Add2~17_sumout\ & \R.aluOp.ALUOpSub~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101000001010000010100000101111111110000010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add2~17_sumout\,
	datac => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datad => \ALT_INV_Selector31~6_OTERM381\,
	dataf => \ALT_INV_ShiftRight1~39_combout\,
	combout => \vAluRes~4_RESYN1068_BDD1069\);

-- Location: LABCELL_X80_Y8_N30
\vAluRes~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~4_combout\ = ( \vAluRes~4_RESYN1068_BDD1069\ & ( \Add1~17_sumout\ & ( (\R.aluRes[4]~DUPLICATE_q\) # (\R.aluCalc~q\) ) ) ) # ( !\vAluRes~4_RESYN1068_BDD1069\ & ( \Add1~17_sumout\ & ( (!\R.aluCalc~q\ & (((\R.aluRes[4]~DUPLICATE_q\)))) # 
-- (\R.aluCalc~q\ & ((!\Selector28~3_combout\) # ((\R.aluOp.ALUOpAdd~q\)))) ) ) ) # ( \vAluRes~4_RESYN1068_BDD1069\ & ( !\Add1~17_sumout\ & ( (\R.aluRes[4]~DUPLICATE_q\) # (\R.aluCalc~q\) ) ) ) # ( !\vAluRes~4_RESYN1068_BDD1069\ & ( !\Add1~17_sumout\ & ( 
-- (!\R.aluCalc~q\ & ((\R.aluRes[4]~DUPLICATE_q\))) # (\R.aluCalc~q\ & (!\Selector28~3_combout\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010111000101110001111110011111100101110001111110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector28~3_combout\,
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_R.aluRes[4]~DUPLICATE_q\,
	datad => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datae => \ALT_INV_vAluRes~4_RESYN1068_BDD1069\,
	dataf => \ALT_INV_Add1~17_sumout\,
	combout => \vAluRes~4_combout\);

-- Location: LABCELL_X80_Y6_N39
\Comb:vJumpAdr[4]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[4]~0_combout\ = ( \Add3~17_sumout\ & ( (!\Equal4~2_combout\) # (\vAluRes~4_combout\) ) ) # ( !\Add3~17_sumout\ & ( (\vAluRes~4_combout\ & \Equal4~2_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101000001010000010111110101111101011111010111110101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluRes~4_combout\,
	datac => \ALT_INV_Equal4~2_combout\,
	dataf => \ALT_INV_Add3~17_sumout\,
	combout => \Comb:vJumpAdr[4]~0_combout\);

-- Location: FF_X80_Y6_N40
\R.curPC[4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[4]~0_combout\,
	asdata => \Add0~9_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(4));

-- Location: LABCELL_X80_Y6_N27
\R.regWriteData[4]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.regWriteData[4]~feeder_combout\ = \Add0~9_sumout\

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101010101010101010101010101010101010101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add0~9_sumout\,
	combout => \R.regWriteData[4]~feeder_combout\);

-- Location: IOIBUF_X89_Y21_N38
\avm_d_readdata[28]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(28),
	o => \avm_d_readdata[28]~input_o\);

-- Location: FF_X80_Y6_N17
\R.aluRes[4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector28~4_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(4));

-- Location: LABCELL_X80_Y6_N18
\Comb:vRegWriteData[4]~0_RESYN1090\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[4]~0_RESYN1090_BDD1091\ = ( \ShiftRight1~39_combout\ & ( \R.aluRes\(4) & ( (!\R.memToReg~q\ & ((!\R.aluCalc~q\) # ((\Selector31~6_OTERM381\)))) # (\R.memToReg~q\ & (((\Mux222~0_combout\)))) ) ) ) # ( !\ShiftRight1~39_combout\ & ( 
-- \R.aluRes\(4) & ( (!\R.memToReg~q\ & (!\R.aluCalc~q\)) # (\R.memToReg~q\ & ((\Mux222~0_combout\))) ) ) ) # ( \ShiftRight1~39_combout\ & ( !\R.aluRes\(4) & ( (!\R.memToReg~q\ & (\R.aluCalc~q\ & ((\Selector31~6_OTERM381\)))) # (\R.memToReg~q\ & 
-- (((\Mux222~0_combout\)))) ) ) ) # ( !\ShiftRight1~39_combout\ & ( !\R.aluRes\(4) & ( (\Mux222~0_combout\ & \R.memToReg~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000110101001110100011101000111010001111110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluCalc~q\,
	datab => \ALT_INV_Mux222~0_combout\,
	datac => \ALT_INV_R.memToReg~q\,
	datad => \ALT_INV_Selector31~6_OTERM381\,
	datae => \ALT_INV_ShiftRight1~39_combout\,
	dataf => \ALT_INV_R.aluRes\(4),
	combout => \Comb:vRegWriteData[4]~0_RESYN1090_BDD1091\);

-- Location: LABCELL_X80_Y6_N42
\Comb:vRegWriteData[4]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[4]~0_combout\ = ( \Selector28~3_combout\ & ( \Comb:vRegWriteData[4]~0_RESYN1090_BDD1091\ & ( (!\R.memToReg~q\) # (\avm_d_readdata[28]~input_o\) ) ) ) # ( !\Selector28~3_combout\ & ( \Comb:vRegWriteData[4]~0_RESYN1090_BDD1091\ & ( 
-- (!\R.memToReg~q\) # (\avm_d_readdata[28]~input_o\) ) ) ) # ( \Selector28~3_combout\ & ( !\Comb:vRegWriteData[4]~0_RESYN1090_BDD1091\ & ( (!\R.memToReg~q\ & (\Selector28~0_combout\ & \R.aluCalc~q\)) ) ) ) # ( !\Selector28~3_combout\ & ( 
-- !\Comb:vRegWriteData[4]~0_RESYN1090_BDD1091\ & ( (!\R.memToReg~q\ & \R.aluCalc~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000010101010000000000000101010111011101110111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.memToReg~q\,
	datab => \ALT_INV_avm_d_readdata[28]~input_o\,
	datac => \ALT_INV_Selector28~0_combout\,
	datad => \ALT_INV_R.aluCalc~q\,
	datae => \ALT_INV_Selector28~3_combout\,
	dataf => \ALT_INV_Comb:vRegWriteData[4]~0_RESYN1090_BDD1091\,
	combout => \Comb:vRegWriteData[4]~0_combout\);

-- Location: FF_X80_Y6_N29
\R.regWriteData[4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \R.regWriteData[4]~feeder_combout\,
	asdata => \Comb:vRegWriteData[4]~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(4));

-- Location: LABCELL_X62_Y7_N18
\RegFile[23][4]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \RegFile[23][4]~feeder_combout\ = ( \R.regWriteData\(4) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_R.regWriteData\(4),
	combout => \RegFile[23][4]~feeder_combout\);

-- Location: FF_X62_Y7_N19
\RegFile[23][4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[23][4]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~12_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[23][4]~q\);

-- Location: LABCELL_X63_Y5_N18
\Mux118~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux118~18_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[16][4]~q\))) # (\R.curInst\(20) & (\RegFile[17][4]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[18][4]~q\))) # (\R.curInst\(20) & (\RegFile[19][4]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[17][4]~q\,
	datab => \ALT_INV_RegFile[19][4]~q\,
	datac => \ALT_INV_RegFile[18][4]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][4]~q\,
	combout => \Mux118~18_combout\);

-- Location: LABCELL_X64_Y5_N48
\Mux118~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux118~5_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux118~18_combout\))))) # (\R.curInst\(22) & (((!\Mux118~18_combout\ & (\RegFile[20][4]~q\)) # (\Mux118~18_combout\ & ((\RegFile[21][4]~q\)))))) ) ) # ( \R.curInst\(21) & ( 
-- (!\R.curInst\(22) & ((((\Mux118~18_combout\))))) # (\R.curInst\(22) & (((!\Mux118~18_combout\ & ((\RegFile[22][4]~q\))) # (\Mux118~18_combout\ & (\RegFile[23][4]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110101010111111111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[23][4]~q\,
	datac => \ALT_INV_RegFile[22][4]~q\,
	datad => \ALT_INV_RegFile[21][4]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux118~18_combout\,
	datag => \ALT_INV_RegFile[20][4]~q\,
	combout => \Mux118~5_combout\);

-- Location: LABCELL_X64_Y5_N42
\Mux118~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux118~14_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[8][4]~q\))) # (\R.curInst\(20) & (\RegFile[9][4]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[10][4]~q\))) # (\R.curInst\(20) & (\RegFile[11][4]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][4]~q\,
	datab => \ALT_INV_RegFile[11][4]~q\,
	datac => \ALT_INV_RegFile[10][4]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][4]~q\,
	combout => \Mux118~14_combout\);

-- Location: LABCELL_X64_Y5_N54
\Mux118~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux118~1_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux118~14_combout\)))) # (\R.curInst\(22) & ((!\Mux118~14_combout\ & ((\RegFile[12][4]~q\))) # (\Mux118~14_combout\ & (\RegFile[13][4]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux118~14_combout\)))) # (\R.curInst\(22) & ((!\Mux118~14_combout\ & ((\RegFile[14][4]~q\))) # (\Mux118~14_combout\ & (\RegFile[15][4]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][4]~q\,
	datab => \ALT_INV_RegFile[13][4]~q\,
	datac => \ALT_INV_RegFile[14][4]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux118~14_combout\,
	datag => \ALT_INV_RegFile[12][4]~q\,
	combout => \Mux118~1_combout\);

-- Location: MLABCELL_X65_Y7_N30
\Mux118~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux118~0_combout\ = ( \RegFile[5][4]~q\ & ( \R.curInst\(21) & ( (!\R.curInst\(20) & (\RegFile[6][4]~q\)) # (\R.curInst\(20) & ((\RegFile[7][4]~q\))) ) ) ) # ( !\RegFile[5][4]~q\ & ( \R.curInst\(21) & ( (!\R.curInst\(20) & (\RegFile[6][4]~q\)) # 
-- (\R.curInst\(20) & ((\RegFile[7][4]~q\))) ) ) ) # ( \RegFile[5][4]~q\ & ( !\R.curInst\(21) & ( (\R.curInst\(20)) # (\RegFile[4][4]~q\) ) ) ) # ( !\RegFile[5][4]~q\ & ( !\R.curInst\(21) & ( (\RegFile[4][4]~q\ & !\R.curInst\(20)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010100000000010101011111111100110011000011110011001100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[4][4]~q\,
	datab => \ALT_INV_RegFile[6][4]~q\,
	datac => \ALT_INV_RegFile[7][4]~q\,
	datad => \ALT_INV_R.curInst\(20),
	datae => \ALT_INV_RegFile[5][4]~q\,
	dataf => \ALT_INV_R.curInst\(21),
	combout => \Mux118~0_combout\);

-- Location: MLABCELL_X65_Y7_N0
\Mux118~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux118~26_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (\RegFile[1][4]~q\ & (\R.curInst\(20)))) # (\R.curInst\(22) & (((\Mux118~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (((\RegFile[2][4]~q\)))) # 
-- (\R.curInst\(20) & (\RegFile[3][4]~q\)))) # (\R.curInst\(22) & ((((\Mux118~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001100000011000100010000110011001111110011111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][4]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[2][4]~q\,
	datad => \ALT_INV_R.curInst\(20),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux118~0_combout\,
	datag => \ALT_INV_RegFile[1][4]~q\,
	combout => \Mux118~26_combout\);

-- Location: LABCELL_X61_Y3_N48
\Mux118~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux118~22_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[24][4]~q\))) # (\R.curInst\(20) & (\RegFile[25][4]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[26][4]~q\))) # (\R.curInst\(20) & (\RegFile[27][4]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[25][4]~q\,
	datab => \ALT_INV_RegFile[27][4]~q\,
	datac => \ALT_INV_RegFile[26][4]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][4]~q\,
	combout => \Mux118~22_combout\);

-- Location: LABCELL_X61_Y3_N42
\Mux118~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux118~9_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux118~22_combout\)))) # (\R.curInst\(22) & ((!\Mux118~22_combout\ & ((\RegFile[28][4]~q\))) # (\Mux118~22_combout\ & (\RegFile[29][4]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux118~22_combout\)))) # (\R.curInst\(22) & ((!\Mux118~22_combout\ & ((\RegFile[30][4]~q\))) # (\Mux118~22_combout\ & (\RegFile[31][4]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][4]~q\,
	datab => \ALT_INV_RegFile[29][4]~q\,
	datac => \ALT_INV_RegFile[30][4]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux118~22_combout\,
	datag => \ALT_INV_RegFile[28][4]~q\,
	combout => \Mux118~9_combout\);

-- Location: LABCELL_X64_Y5_N18
\Mux118~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux118~13_combout\ = ( \Mux118~26_combout\ & ( \Mux118~9_combout\ & ( (!\R.curInst\(23) & (((!\R.curInst\(24))) # (\Mux118~5_combout\))) # (\R.curInst\(23) & (((\R.curInst\(24)) # (\Mux118~1_combout\)))) ) ) ) # ( !\Mux118~26_combout\ & ( 
-- \Mux118~9_combout\ & ( (!\R.curInst\(23) & (\Mux118~5_combout\ & ((\R.curInst\(24))))) # (\R.curInst\(23) & (((\R.curInst\(24)) # (\Mux118~1_combout\)))) ) ) ) # ( \Mux118~26_combout\ & ( !\Mux118~9_combout\ & ( (!\R.curInst\(23) & (((!\R.curInst\(24))) # 
-- (\Mux118~5_combout\))) # (\R.curInst\(23) & (((\Mux118~1_combout\ & !\R.curInst\(24))))) ) ) ) # ( !\Mux118~26_combout\ & ( !\Mux118~9_combout\ & ( (!\R.curInst\(23) & (\Mux118~5_combout\ & ((\R.curInst\(24))))) # (\R.curInst\(23) & (((\Mux118~1_combout\ 
-- & !\R.curInst\(24))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001101000100110011110100010000000011011101111100111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux118~5_combout\,
	datab => \ALT_INV_R.curInst\(23),
	datac => \ALT_INV_Mux118~1_combout\,
	datad => \ALT_INV_R.curInst\(24),
	datae => \ALT_INV_Mux118~26_combout\,
	dataf => \ALT_INV_Mux118~9_combout\,
	combout => \Mux118~13_combout\);

-- Location: MLABCELL_X72_Y5_N27
\NxR.aluData2[4]~20\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[4]~20_combout\ = ( \Mux118~13_combout\ & ( (!\vAluSrc2~1_combout\) # ((\Equal4~1_combout\ & \Mux150~0_combout\)) ) ) # ( !\Mux118~13_combout\ & ( (\vAluSrc2~1_combout\ & (\Equal4~1_combout\ & \Mux150~0_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000100000001000000010000000110101011101010111010101110101011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluSrc2~1_combout\,
	datab => \ALT_INV_Equal4~1_combout\,
	datac => \ALT_INV_Mux150~0_combout\,
	dataf => \ALT_INV_Mux118~13_combout\,
	combout => \NxR.aluData2[4]~20_combout\);

-- Location: LABCELL_X71_Y9_N12
\Selector12~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector12~2_combout\ = ( \R.aluOp.ALUOpSLL_OTERM359\ & ( \NxR.aluData2[4]~20_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000001111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datae => \ALT_INV_R.aluOp.ALUOpSLL_OTERM359\,
	dataf => \ALT_INV_NxR.aluData2[4]~20_combout\,
	combout => \Selector12~2_combout\);

-- Location: FF_X71_Y9_N13
\Selector12~2_NEW_REG394\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector12~2_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector12~2_OTERM395\);

-- Location: LABCELL_X81_Y7_N12
\Selector11~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector11~2_combout\ = ( \R.aluData1\(21) & ( \R.aluOp.ALUOpXor~DUPLICATE_q\ & ( (!\R.aluData2\(21)) # ((\R.aluData2\(4) & (\R.aluData1\(31) & \R.aluOp.ALUOpSRA~q\))) ) ) ) # ( !\R.aluData1\(21) & ( \R.aluOp.ALUOpXor~DUPLICATE_q\ & ( ((\R.aluData2\(4) & 
-- (\R.aluData1\(31) & \R.aluOp.ALUOpSRA~q\))) # (\R.aluData2\(21)) ) ) ) # ( \R.aluData1\(21) & ( !\R.aluOp.ALUOpXor~DUPLICATE_q\ & ( (\R.aluData2\(4) & (\R.aluData1\(31) & \R.aluOp.ALUOpSRA~q\)) ) ) ) # ( !\R.aluData1\(21) & ( 
-- !\R.aluOp.ALUOpXor~DUPLICATE_q\ & ( (\R.aluData2\(4) & (\R.aluData1\(31) & \R.aluOp.ALUOpSRA~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000011000000000000001101010101010101111010101010101011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(21),
	datab => \ALT_INV_R.aluData2\(4),
	datac => \ALT_INV_R.aluData1\(31),
	datad => \ALT_INV_R.aluOp.ALUOpSRA~q\,
	datae => \ALT_INV_R.aluData1\(21),
	dataf => \ALT_INV_R.aluOp.ALUOpXor~DUPLICATE_q\,
	combout => \Selector11~2_combout\);

-- Location: MLABCELL_X84_Y7_N57
\Selector11~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector11~3_combout\ = ( \R.aluData2\(21) & ( \R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( (\R.aluOp.ALUOpOr~q\) # (\R.aluData1\(21)) ) ) ) # ( !\R.aluData2\(21) & ( \R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( (\R.aluData1\(21) & \R.aluOp.ALUOpOr~q\) ) ) ) # ( 
-- \R.aluData2\(21) & ( !\R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( \R.aluOp.ALUOpOr~q\ ) ) ) # ( !\R.aluData2\(21) & ( !\R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( (\R.aluData1\(21) & \R.aluOp.ALUOpOr~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101000011110000111100000101000001010101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData1\(21),
	datac => \ALT_INV_R.aluOp.ALUOpOr~q\,
	datae => \ALT_INV_R.aluData2\(21),
	dataf => \ALT_INV_R.aluOp.ALUOpAnd~DUPLICATE_q\,
	combout => \Selector11~3_combout\);

-- Location: LABCELL_X81_Y7_N54
\Selector11~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector11~4_combout\ = ( \ShiftLeft0~6_OTERM243\ & ( !\Selector11~3_combout\ & ( (!\Selector12~2_OTERM395\ & !\Selector11~2_combout\) ) ) ) # ( !\ShiftLeft0~6_OTERM243\ & ( !\Selector11~3_combout\ & ( (!\Selector11~2_combout\ & 
-- ((!\Selector12~2_OTERM395\) # ((!\ShiftLeft0~7_OTERM205\) # (\ShiftRight0~7_OTERM233DUPLICATE_q\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1100100011001100100010001000100000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector12~2_OTERM395\,
	datab => \ALT_INV_Selector11~2_combout\,
	datac => \ALT_INV_ShiftLeft0~7_OTERM205\,
	datad => \ALT_INV_ShiftRight0~7_OTERM233DUPLICATE_q\,
	datae => \ALT_INV_ShiftLeft0~6_OTERM243\,
	dataf => \ALT_INV_Selector11~3_combout\,
	combout => \Selector11~4_combout\);

-- Location: MLABCELL_X78_Y2_N54
\Selector11~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector11~5_combout\ = ( \R.aluOp.ALUOpAdd~q\ & ( \Add2~85_sumout\ & ( (!\Selector11~4_combout\) # (((\Add1~85_sumout\) # (\Selector11~1_combout\)) # (\R.aluOp.ALUOpSub~q\)) ) ) ) # ( !\R.aluOp.ALUOpAdd~q\ & ( \Add2~85_sumout\ & ( 
-- (!\Selector11~4_combout\) # ((\Selector11~1_combout\) # (\R.aluOp.ALUOpSub~q\)) ) ) ) # ( \R.aluOp.ALUOpAdd~q\ & ( !\Add2~85_sumout\ & ( (!\Selector11~4_combout\) # ((\Add1~85_sumout\) # (\Selector11~1_combout\)) ) ) ) # ( !\R.aluOp.ALUOpAdd~q\ & ( 
-- !\Add2~85_sumout\ & ( (!\Selector11~4_combout\) # (\Selector11~1_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010111110101111101011111111111110111111101111111011111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector11~4_combout\,
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_Selector11~1_combout\,
	datad => \ALT_INV_Add1~85_sumout\,
	datae => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	dataf => \ALT_INV_Add2~85_sumout\,
	combout => \Selector11~5_combout\);

-- Location: MLABCELL_X78_Y2_N33
\Comb:vJumpAdr[21]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[21]~0_combout\ = ( \R.aluRes\(21) & ( \Add3~85_sumout\ & ( (!\R.aluCalc~q\) # ((!\Equal4~2_combout\) # (\Selector11~5_combout\)) ) ) ) # ( !\R.aluRes\(21) & ( \Add3~85_sumout\ & ( (!\Equal4~2_combout\) # ((\R.aluCalc~q\ & 
-- \Selector11~5_combout\)) ) ) ) # ( \R.aluRes\(21) & ( !\Add3~85_sumout\ & ( (\Equal4~2_combout\ & ((!\R.aluCalc~q\) # (\Selector11~5_combout\))) ) ) ) # ( !\R.aluRes\(21) & ( !\Add3~85_sumout\ & ( (\R.aluCalc~q\ & (\Selector11~5_combout\ & 
-- \Equal4~2_combout\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000100000001000010110000101111110001111100011111101111111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluCalc~q\,
	datab => \ALT_INV_Selector11~5_combout\,
	datac => \ALT_INV_Equal4~2_combout\,
	datae => \ALT_INV_R.aluRes\(21),
	dataf => \ALT_INV_Add3~85_sumout\,
	combout => \Comb:vJumpAdr[21]~0_combout\);

-- Location: FF_X78_Y2_N34
\R.curPC[21]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[21]~0_combout\,
	asdata => \Add0~77_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC[21]~DUPLICATE_q\);

-- Location: MLABCELL_X78_Y2_N39
\R.regWriteData[21]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.regWriteData[21]~feeder_combout\ = ( \Add0~77_sumout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \ALT_INV_Add0~77_sumout\,
	combout => \R.regWriteData[21]~feeder_combout\);

-- Location: LABCELL_X80_Y4_N21
\Comb:vRegWriteData[21]~1_RESYN1130\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[21]~1_RESYN1130_BDD1131\ = (\R.aluCalc~q\ & !\R.memToReg~q\)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100000000001100110000000000110011000000000011001100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluCalc~q\,
	datad => \ALT_INV_R.memToReg~q\,
	combout => \Comb:vRegWriteData[21]~1_RESYN1130_BDD1131\);

-- Location: IOIBUF_X84_Y0_N1
\avm_d_readdata[13]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(13),
	o => \avm_d_readdata[13]~input_o\);

-- Location: LABCELL_X79_Y2_N6
\Comb:vRegWriteData[21]~1_RESYN1126\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[21]~1_RESYN1126_BDD1127\ = ( \avm_d_readdata[23]~input_o\ & ( \avm_d_readdata[13]~input_o\ & ( (!\R.curInst\(14) & ((!\R.curInst\(12) & ((\R.curInst\(13)) # (\avm_d_readdata[31]~input_o\))) # (\R.curInst\(12) & ((!\R.curInst\(13)))))) 
-- ) ) ) # ( !\avm_d_readdata[23]~input_o\ & ( \avm_d_readdata[13]~input_o\ & ( (!\R.curInst\(12) & (!\R.curInst\(14) & ((\R.curInst\(13)) # (\avm_d_readdata[31]~input_o\)))) ) ) ) # ( \avm_d_readdata[23]~input_o\ & ( !\avm_d_readdata[13]~input_o\ & ( 
-- (!\R.curInst\(13) & (!\R.curInst\(14) & ((\avm_d_readdata[31]~input_o\) # (\R.curInst\(12))))) ) ) ) # ( !\avm_d_readdata[23]~input_o\ & ( !\avm_d_readdata[13]~input_o\ & ( (!\R.curInst\(12) & (\avm_d_readdata[31]~input_o\ & (!\R.curInst\(13) & 
-- !\R.curInst\(14)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010000000000000011100000000000000101010000000000111101000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(12),
	datab => \ALT_INV_avm_d_readdata[31]~input_o\,
	datac => \ALT_INV_R.curInst\(13),
	datad => \ALT_INV_R.curInst\(14),
	datae => \ALT_INV_avm_d_readdata[23]~input_o\,
	dataf => \ALT_INV_avm_d_readdata[13]~input_o\,
	combout => \Comb:vRegWriteData[21]~1_RESYN1126_BDD1127\);

-- Location: MLABCELL_X78_Y2_N24
\Comb:vRegWriteData[21]~1_RESYN1128\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[21]~1_RESYN1128_BDD1129\ = ( \Comb:vRegWriteData[21]~1_RESYN1126_BDD1127\ & ( \Add2~85_sumout\ & ( ((!\R.aluCalc~q\ & ((\R.aluRes\(21)))) # (\R.aluCalc~q\ & (\R.aluOp.ALUOpSub~q\))) # (\R.memToReg~q\) ) ) ) # ( 
-- !\Comb:vRegWriteData[21]~1_RESYN1126_BDD1127\ & ( \Add2~85_sumout\ & ( (!\R.memToReg~q\ & ((!\R.aluCalc~q\ & ((\R.aluRes\(21)))) # (\R.aluCalc~q\ & (\R.aluOp.ALUOpSub~q\)))) ) ) ) # ( \Comb:vRegWriteData[21]~1_RESYN1126_BDD1127\ & ( !\Add2~85_sumout\ & ( 
-- ((\R.aluRes\(21) & !\R.aluCalc~q\)) # (\R.memToReg~q\) ) ) ) # ( !\Comb:vRegWriteData[21]~1_RESYN1126_BDD1127\ & ( !\Add2~85_sumout\ & ( (!\R.memToReg~q\ & (\R.aluRes\(21) & !\R.aluCalc~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101000000000010111110101010100001010001000100101111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.memToReg~q\,
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_R.aluRes\(21),
	datad => \ALT_INV_R.aluCalc~q\,
	datae => \ALT_INV_Comb:vRegWriteData[21]~1_RESYN1126_BDD1127\,
	dataf => \ALT_INV_Add2~85_sumout\,
	combout => \Comb:vRegWriteData[21]~1_RESYN1128_BDD1129\);

-- Location: MLABCELL_X78_Y2_N48
\Comb:vRegWriteData[21]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[21]~1_combout\ = ( \Selector11~1_combout\ & ( \Comb:vRegWriteData[21]~1_RESYN1128_BDD1129\ ) ) # ( !\Selector11~1_combout\ & ( \Comb:vRegWriteData[21]~1_RESYN1128_BDD1129\ ) ) # ( \Selector11~1_combout\ & ( 
-- !\Comb:vRegWriteData[21]~1_RESYN1128_BDD1129\ & ( \Comb:vRegWriteData[21]~1_RESYN1130_BDD1131\ ) ) ) # ( !\Selector11~1_combout\ & ( !\Comb:vRegWriteData[21]~1_RESYN1128_BDD1129\ & ( (\Comb:vRegWriteData[21]~1_RESYN1130_BDD1131\ & 
-- ((!\Selector11~4_combout\) # ((\R.aluOp.ALUOpAdd~q\ & \Add1~85_sumout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101000001010001010101010101010111111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Comb:vRegWriteData[21]~1_RESYN1130_BDD1131\,
	datab => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datac => \ALT_INV_Selector11~4_combout\,
	datad => \ALT_INV_Add1~85_sumout\,
	datae => \ALT_INV_Selector11~1_combout\,
	dataf => \ALT_INV_Comb:vRegWriteData[21]~1_RESYN1128_BDD1129\,
	combout => \Comb:vRegWriteData[21]~1_combout\);

-- Location: FF_X78_Y2_N41
\R.regWriteData[21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \R.regWriteData[21]~feeder_combout\,
	asdata => \Comb:vRegWriteData[21]~1_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(21));

-- Location: FF_X62_Y3_N38
\RegFile[3][21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(21),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][21]~q\);

-- Location: LABCELL_X62_Y3_N48
\Mux101~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux101~0_combout\ = ( \RegFile[5][21]~q\ & ( \R.curInst\(21) & ( (!\R.curInst\(20) & ((\RegFile[6][21]~q\))) # (\R.curInst\(20) & (\RegFile[7][21]~q\)) ) ) ) # ( !\RegFile[5][21]~q\ & ( \R.curInst\(21) & ( (!\R.curInst\(20) & ((\RegFile[6][21]~q\))) # 
-- (\R.curInst\(20) & (\RegFile[7][21]~q\)) ) ) ) # ( \RegFile[5][21]~q\ & ( !\R.curInst\(21) & ( (\RegFile[4][21]~q\) # (\R.curInst\(20)) ) ) ) # ( !\RegFile[5][21]~q\ & ( !\R.curInst\(21) & ( (!\R.curInst\(20) & \RegFile[4][21]~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101000001010010111110101111100010001101110110001000110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(20),
	datab => \ALT_INV_RegFile[7][21]~q\,
	datac => \ALT_INV_RegFile[4][21]~q\,
	datad => \ALT_INV_RegFile[6][21]~q\,
	datae => \ALT_INV_RegFile[5][21]~q\,
	dataf => \ALT_INV_R.curInst\(21),
	combout => \Mux101~0_combout\);

-- Location: LABCELL_X61_Y5_N0
\Mux101~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux101~26_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((\RegFile[1][21]~q\ & (\R.curInst\(20)))))) # (\R.curInst\(22) & ((((\Mux101~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (((\RegFile[2][21]~q\)))) 
-- # (\R.curInst\(20) & (\RegFile[3][21]~q\)))) # (\R.curInst\(22) & ((((\Mux101~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001010000010100010001001010101010111110101111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[3][21]~q\,
	datac => \ALT_INV_RegFile[2][21]~q\,
	datad => \ALT_INV_R.curInst\(20),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux101~0_combout\,
	datag => \ALT_INV_RegFile[1][21]~q\,
	combout => \Mux101~26_combout\);

-- Location: LABCELL_X64_Y3_N36
\Mux101~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux101~14_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[8][21]~q\))) # (\R.curInst\(20) & (\RegFile[9][21]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[10][21]~q\))) # (\R.curInst\(20) & (\RegFile[11][21]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000001010101111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][21]~q\,
	datab => \ALT_INV_RegFile[11][21]~q\,
	datac => \ALT_INV_RegFile[10][21]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][21]~q\,
	combout => \Mux101~14_combout\);

-- Location: MLABCELL_X65_Y5_N0
\Mux101~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux101~1_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux101~14_combout\)))) # (\R.curInst\(22) & ((!\Mux101~14_combout\ & ((\RegFile[12][21]~q\))) # (\Mux101~14_combout\ & (\RegFile[13][21]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux101~14_combout\)))) # (\R.curInst\(22) & ((!\Mux101~14_combout\ & ((\RegFile[14][21]~q\))) # (\Mux101~14_combout\ & (\RegFile[15][21]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][21]~q\,
	datab => \ALT_INV_RegFile[15][21]~q\,
	datac => \ALT_INV_RegFile[14][21]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux101~14_combout\,
	datag => \ALT_INV_RegFile[12][21]~q\,
	combout => \Mux101~1_combout\);

-- Location: LABCELL_X64_Y1_N12
\Mux101~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux101~18_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & (\RegFile[16][21]~q\)) # (\R.curInst\(20) & ((\RegFile[17][21]~q\)))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & ((\RegFile[18][21]~q\))) # (\R.curInst\(20) & (\RegFile[19][21]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001010101111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[19][21]~q\,
	datac => \ALT_INV_RegFile[18][21]~q\,
	datad => \ALT_INV_RegFile[17][21]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][21]~q\,
	combout => \Mux101~18_combout\);

-- Location: LABCELL_X62_Y5_N12
\Mux101~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux101~5_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux101~18_combout\)))) # (\R.curInst\(22) & ((!\Mux101~18_combout\ & ((\RegFile[20][21]~q\))) # (\Mux101~18_combout\ & (\RegFile[21][21]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux101~18_combout\)))) # (\R.curInst\(22) & ((!\Mux101~18_combout\ & ((\RegFile[22][21]~q\))) # (\Mux101~18_combout\ & (\RegFile[23][21]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[23][21]~q\,
	datab => \ALT_INV_RegFile[21][21]~q\,
	datac => \ALT_INV_RegFile[22][21]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux101~18_combout\,
	datag => \ALT_INV_RegFile[20][21]~q\,
	combout => \Mux101~5_combout\);

-- Location: LABCELL_X62_Y2_N48
\Mux101~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux101~22_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[24][21]~q\))) # (\R.curInst\(20) & (\RegFile[25][21]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & (\RegFile[26][21]~q\)) # (\R.curInst\(20) & ((\RegFile[27][21]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[25][21]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[26][21]~q\,
	datad => \ALT_INV_RegFile[27][21]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][21]~q\,
	combout => \Mux101~22_combout\);

-- Location: LABCELL_X62_Y5_N30
\Mux101~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux101~9_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux101~22_combout\)))) # (\R.curInst\(22) & ((!\Mux101~22_combout\ & ((\RegFile[28][21]~q\))) # (\Mux101~22_combout\ & (\RegFile[29][21]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux101~22_combout\)))) # (\R.curInst\(22) & ((!\Mux101~22_combout\ & ((\RegFile[30][21]~q\))) # (\Mux101~22_combout\ & (\RegFile[31][21]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][21]~q\,
	datab => \ALT_INV_RegFile[29][21]~q\,
	datac => \ALT_INV_RegFile[30][21]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux101~22_combout\,
	datag => \ALT_INV_RegFile[28][21]~q\,
	combout => \Mux101~9_combout\);

-- Location: LABCELL_X61_Y5_N24
\Mux101~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux101~13_combout\ = ( \Mux101~5_combout\ & ( \Mux101~9_combout\ & ( ((!\R.curInst\(23) & (\Mux101~26_combout\)) # (\R.curInst\(23) & ((\Mux101~1_combout\)))) # (\R.curInst\(24)) ) ) ) # ( !\Mux101~5_combout\ & ( \Mux101~9_combout\ & ( (!\R.curInst\(23) 
-- & (\Mux101~26_combout\ & ((!\R.curInst\(24))))) # (\R.curInst\(23) & (((\R.curInst\(24)) # (\Mux101~1_combout\)))) ) ) ) # ( \Mux101~5_combout\ & ( !\Mux101~9_combout\ & ( (!\R.curInst\(23) & (((\R.curInst\(24))) # (\Mux101~26_combout\))) # 
-- (\R.curInst\(23) & (((\Mux101~1_combout\ & !\R.curInst\(24))))) ) ) ) # ( !\Mux101~5_combout\ & ( !\Mux101~9_combout\ & ( (!\R.curInst\(24) & ((!\R.curInst\(23) & (\Mux101~26_combout\)) # (\R.curInst\(23) & ((\Mux101~1_combout\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100011100000000010001111100110001000111001100110100011111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux101~26_combout\,
	datab => \ALT_INV_R.curInst\(23),
	datac => \ALT_INV_Mux101~1_combout\,
	datad => \ALT_INV_R.curInst\(24),
	datae => \ALT_INV_Mux101~5_combout\,
	dataf => \ALT_INV_Mux101~9_combout\,
	combout => \Mux101~13_combout\);

-- Location: LABCELL_X74_Y5_N54
\NxR.aluData2[21]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[21]~0_combout\ = ( \Mux133~0_combout\ & ( (!\vAluSrc2~1_combout\ & ((\Mux101~13_combout\))) # (\vAluSrc2~1_combout\ & (\Equal4~1_combout\)) ) ) # ( !\Mux133~0_combout\ & ( (!\vAluSrc2~1_combout\ & \Mux101~13_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011110000000000001111000000000011111100110000001111110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Equal4~1_combout\,
	datac => \ALT_INV_vAluSrc2~1_combout\,
	datad => \ALT_INV_Mux101~13_combout\,
	dataf => \ALT_INV_Mux133~0_combout\,
	combout => \NxR.aluData2[21]~0_combout\);

-- Location: FF_X74_Y5_N10
\R.aluData2[21]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \NxR.aluData2[21]~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData2\(21));

-- Location: MLABCELL_X78_Y5_N6
\Add1~89\ : cyclonev_lcell_comb
-- Equation(s):
-- \Add1~89_sumout\ = SUM(( \R.aluData2\(22) ) + ( \R.aluData1\(22) ) + ( \Add1~86\ ))
-- \Add1~90\ = CARRY(( \R.aluData2\(22) ) + ( \R.aluData1\(22) ) + ( \Add1~86\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluData2\(22),
	datac => \ALT_INV_R.aluData1\(22),
	cin => \Add1~86\,
	sumout => \Add1~89_sumout\,
	cout => \Add1~90\);

-- Location: LABCELL_X77_Y2_N42
\Comb:vJumpAdr[22]~0_RESYN1028\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[22]~0_RESYN1028_BDD1029\ = ( \Add2~89_sumout\ & ( \Selector10~4_combout\ & ( (!\R.aluCalc~q\ & (\R.aluRes\(22))) # (\R.aluCalc~q\ & (((\Selector10~1_combout\) # (\R.aluOp.ALUOpSub~q\)))) ) ) ) # ( !\Add2~89_sumout\ & ( 
-- \Selector10~4_combout\ & ( (!\R.aluCalc~q\ & (\R.aluRes\(22))) # (\R.aluCalc~q\ & ((\Selector10~1_combout\))) ) ) ) # ( \Add2~89_sumout\ & ( !\Selector10~4_combout\ & ( (\R.aluCalc~q\) # (\R.aluRes\(22)) ) ) ) # ( !\Add2~89_sumout\ & ( 
-- !\Selector10~4_combout\ & ( (\R.aluCalc~q\) # (\R.aluRes\(22)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0111011101110111011101110111011101000100011101110100011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluRes\(22),
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datad => \ALT_INV_Selector10~1_combout\,
	datae => \ALT_INV_Add2~89_sumout\,
	dataf => \ALT_INV_Selector10~4_combout\,
	combout => \Comb:vJumpAdr[22]~0_RESYN1028_BDD1029\);

-- Location: LABCELL_X77_Y2_N12
\Comb:vJumpAdr[22]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[22]~0_combout\ = ( \R.aluOp.ALUOpAdd~q\ & ( \Add3~89_sumout\ & ( (!\Equal4~2_combout\) # (((\R.aluCalc~q\ & \Add1~89_sumout\)) # (\Comb:vJumpAdr[22]~0_RESYN1028_BDD1029\)) ) ) ) # ( !\R.aluOp.ALUOpAdd~q\ & ( \Add3~89_sumout\ & ( 
-- (!\Equal4~2_combout\) # (\Comb:vJumpAdr[22]~0_RESYN1028_BDD1029\) ) ) ) # ( \R.aluOp.ALUOpAdd~q\ & ( !\Add3~89_sumout\ & ( (\Equal4~2_combout\ & (((\R.aluCalc~q\ & \Add1~89_sumout\)) # (\Comb:vJumpAdr[22]~0_RESYN1028_BDD1029\))) ) ) ) # ( 
-- !\R.aluOp.ALUOpAdd~q\ & ( !\Add3~89_sumout\ & ( (\Equal4~2_combout\ & \Comb:vJumpAdr[22]~0_RESYN1028_BDD1029\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110011000000010011001111001100111111111100110111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluCalc~q\,
	datab => \ALT_INV_Equal4~2_combout\,
	datac => \ALT_INV_Add1~89_sumout\,
	datad => \ALT_INV_Comb:vJumpAdr[22]~0_RESYN1028_BDD1029\,
	datae => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	dataf => \ALT_INV_Add3~89_sumout\,
	combout => \Comb:vJumpAdr[22]~0_combout\);

-- Location: FF_X77_Y2_N13
\R.curPC[22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[22]~0_combout\,
	asdata => \Add0~81_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(22));

-- Location: LABCELL_X77_Y2_N24
\Comb:vRegWriteData[22]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[22]~3_combout\ = ( \R.aluCalc~q\ & ( \Selector10~4_combout\ & ( !\Selector10~1_combout\ ) ) ) # ( !\R.aluCalc~q\ & ( \Selector10~4_combout\ & ( (!\R.aluRes\(22) & !\R.memToReg~q\) ) ) ) # ( !\R.aluCalc~q\ & ( !\Selector10~4_combout\ & 
-- ( (!\R.aluRes\(22) & !\R.memToReg~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010000010100000000000000000000010100000101000001100110011001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluRes\(22),
	datab => \ALT_INV_Selector10~1_combout\,
	datac => \ALT_INV_R.memToReg~q\,
	datae => \ALT_INV_R.aluCalc~q\,
	dataf => \ALT_INV_Selector10~4_combout\,
	combout => \Comb:vRegWriteData[22]~3_combout\);

-- Location: IOIBUF_X34_Y0_N58
\avm_d_readdata[14]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(14),
	o => \avm_d_readdata[14]~input_o\);

-- Location: LABCELL_X79_Y1_N27
\Comb:vRegWriteData[22]~2_RESYN1112\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[22]~2_RESYN1112_BDD1113\ = ( \R.curInst\(12) & ( !\avm_d_readdata[23]~input_o\ ) ) # ( !\R.curInst\(12) & ( !\avm_d_readdata[31]~input_o\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1100110011001100110011001100110010101010101010101010101010101010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_avm_d_readdata[23]~input_o\,
	datab => \ALT_INV_avm_d_readdata[31]~input_o\,
	dataf => \ALT_INV_R.curInst\(12),
	combout => \Comb:vRegWriteData[22]~2_RESYN1112_BDD1113\);

-- Location: LABCELL_X79_Y1_N0
\Comb:vRegWriteData[22]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[22]~2_combout\ = ( \Comb:vRegWriteData[22]~2_RESYN1112_BDD1113\ & ( \R.curInst\(12) & ( \R.memToReg~q\ ) ) ) # ( !\Comb:vRegWriteData[22]~2_RESYN1112_BDD1113\ & ( \R.curInst\(12) & ( (\R.memToReg~q\ & ((\R.curInst\(14)) # 
-- (\R.curInst\(13)))) ) ) ) # ( \Comb:vRegWriteData[22]~2_RESYN1112_BDD1113\ & ( !\R.curInst\(12) & ( (\R.memToReg~q\ & ((!\avm_d_readdata[14]~input_o\) # ((!\R.curInst\(13)) # (\R.curInst\(14))))) ) ) ) # ( !\Comb:vRegWriteData[22]~2_RESYN1112_BDD1113\ & ( 
-- !\R.curInst\(12) & ( (\R.memToReg~q\ & (((!\avm_d_readdata[14]~input_o\ & \R.curInst\(13))) # (\R.curInst\(14)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000101111000000001110111100000000001111110000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_avm_d_readdata[14]~input_o\,
	datab => \ALT_INV_R.curInst\(13),
	datac => \ALT_INV_R.curInst\(14),
	datad => \ALT_INV_R.memToReg~q\,
	datae => \ALT_INV_Comb:vRegWriteData[22]~2_RESYN1112_BDD1113\,
	dataf => \ALT_INV_R.curInst\(12),
	combout => \Comb:vRegWriteData[22]~2_combout\);

-- Location: LABCELL_X77_Y2_N18
\Comb:vRegWriteData[22]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[22]~1_combout\ = ( \R.curInst\(13) & ( \Add1~89_sumout\ & ( (!\R.memToReg~q\ & (((\R.aluOp.ALUOpAdd~q\)))) # (\R.memToReg~q\ & (\avm_d_readdata[14]~input_o\ & (!\R.curInst\(14)))) ) ) ) # ( !\R.curInst\(13) & ( \Add1~89_sumout\ & ( 
-- (!\R.memToReg~q\ & ((\R.aluOp.ALUOpAdd~q\))) # (\R.memToReg~q\ & (!\R.curInst\(14))) ) ) ) # ( \R.curInst\(13) & ( !\Add1~89_sumout\ & ( (\avm_d_readdata[14]~input_o\ & (!\R.curInst\(14) & \R.memToReg~q\)) ) ) ) # ( !\R.curInst\(13) & ( !\Add1~89_sumout\ 
-- & ( (!\R.curInst\(14) & \R.memToReg~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000110000001100000001000000010000001100111111000000010011110100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_avm_d_readdata[14]~input_o\,
	datab => \ALT_INV_R.curInst\(14),
	datac => \ALT_INV_R.memToReg~q\,
	datad => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datae => \ALT_INV_R.curInst\(13),
	dataf => \ALT_INV_Add1~89_sumout\,
	combout => \Comb:vRegWriteData[22]~1_combout\);

-- Location: MLABCELL_X78_Y2_N42
\Comb:vRegWriteData[22]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[22]~0_combout\ = ( !\Comb:vRegWriteData[22]~2_combout\ & ( \Comb:vRegWriteData[22]~1_combout\ & ( (!\Comb:vRegWriteData[22]~3_combout\) # (\R.aluCalc~q\) ) ) ) # ( !\Comb:vRegWriteData[22]~2_combout\ & ( 
-- !\Comb:vRegWriteData[22]~1_combout\ & ( (!\Comb:vRegWriteData[22]~3_combout\) # ((\Add2~89_sumout\ & (\R.aluOp.ALUOpSub~q\ & \R.aluCalc~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111100000001000000000000000011111111000011110000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add2~89_sumout\,
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_R.aluCalc~q\,
	datad => \ALT_INV_Comb:vRegWriteData[22]~3_combout\,
	datae => \ALT_INV_Comb:vRegWriteData[22]~2_combout\,
	dataf => \ALT_INV_Comb:vRegWriteData[22]~1_combout\,
	combout => \Comb:vRegWriteData[22]~0_combout\);

-- Location: FF_X81_Y5_N32
\R.regWriteData[22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Add0~81_sumout\,
	asdata => \Comb:vRegWriteData[22]~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(22));

-- Location: FF_X70_Y3_N32
\RegFile[31][22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(22),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~16_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[31][22]~q\);

-- Location: LABCELL_X63_Y2_N18
\Mux100~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux100~22_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[24][22]~q\))) # (\R.curInst\(20) & (\RegFile[25][22]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[26][22]~q\))) # (\R.curInst\(20) & (\RegFile[27][22]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[27][22]~q\,
	datab => \ALT_INV_RegFile[25][22]~q\,
	datac => \ALT_INV_RegFile[26][22]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][22]~q\,
	combout => \Mux100~22_combout\);

-- Location: LABCELL_X63_Y2_N24
\Mux100~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux100~9_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux100~22_combout\)))) # (\R.curInst\(22) & ((!\Mux100~22_combout\ & (\RegFile[28][22]~q\)) # (\Mux100~22_combout\ & ((\RegFile[29][22]~q\)))))) ) ) # ( \R.curInst\(21) & ( 
-- (!\R.curInst\(22) & ((((\Mux100~22_combout\))))) # (\R.curInst\(22) & (((!\Mux100~22_combout\ & ((\RegFile[30][22]~q\))) # (\Mux100~22_combout\ & (\RegFile[31][22]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111001100111111111101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][22]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[30][22]~q\,
	datad => \ALT_INV_RegFile[29][22]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux100~22_combout\,
	datag => \ALT_INV_RegFile[28][22]~q\,
	combout => \Mux100~9_combout\);

-- Location: LABCELL_X68_Y2_N12
\Mux100~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux100~14_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & (\RegFile[8][22]~q\)) # (\R.curInst\(20) & ((\RegFile[9][22]~q\)))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & ((\RegFile[10][22]~q\))) # (\R.curInst\(20) & (\RegFile[11][22]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001010101111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[11][22]~q\,
	datac => \ALT_INV_RegFile[10][22]~q\,
	datad => \ALT_INV_RegFile[9][22]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][22]~q\,
	combout => \Mux100~14_combout\);

-- Location: LABCELL_X62_Y2_N0
\Mux100~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux100~1_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux100~14_combout\)))) # (\R.curInst\(22) & ((!\Mux100~14_combout\ & ((\RegFile[12][22]~q\))) # (\Mux100~14_combout\ & (\RegFile[13][22]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux100~14_combout\)))) # (\R.curInst\(22) & ((!\Mux100~14_combout\ & ((\RegFile[14][22]~q\))) # (\Mux100~14_combout\ & (\RegFile[15][22]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[13][22]~q\,
	datab => \ALT_INV_RegFile[15][22]~q\,
	datac => \ALT_INV_RegFile[14][22]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux100~14_combout\,
	datag => \ALT_INV_RegFile[12][22]~q\,
	combout => \Mux100~1_combout\);

-- Location: LABCELL_X64_Y1_N6
\Mux100~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux100~18_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & (\RegFile[16][22]~q\)) # (\R.curInst\(20) & ((\RegFile[17][22]~q\)))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & ((\RegFile[18][22]~q\))) # (\R.curInst\(20) & (\RegFile[19][22]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001010101111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[19][22]~q\,
	datac => \ALT_INV_RegFile[18][22]~q\,
	datad => \ALT_INV_RegFile[17][22]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][22]~q\,
	combout => \Mux100~18_combout\);

-- Location: LABCELL_X64_Y1_N42
\Mux100~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux100~5_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux100~18_combout\))))) # (\R.curInst\(22) & (((!\Mux100~18_combout\ & ((\RegFile[20][22]~q\))) # (\Mux100~18_combout\ & (\RegFile[21][22]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- (!\R.curInst\(22) & ((((\Mux100~18_combout\))))) # (\R.curInst\(22) & (((!\Mux100~18_combout\ & (\RegFile[22][22]~q\)) # (\Mux100~18_combout\ & ((\RegFile[23][22]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000101000001010000010110111011101110111010101011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[21][22]~q\,
	datac => \ALT_INV_RegFile[22][22]~q\,
	datad => \ALT_INV_RegFile[23][22]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux100~18_combout\,
	datag => \ALT_INV_RegFile[20][22]~q\,
	combout => \Mux100~5_combout\);

-- Location: LABCELL_X68_Y3_N36
\Mux100~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux100~0_combout\ = ( \RegFile[5][22]~q\ & ( \R.curInst\(20) & ( (!\R.curInst\(21)) # (\RegFile[7][22]~q\) ) ) ) # ( !\RegFile[5][22]~q\ & ( \R.curInst\(20) & ( (\R.curInst\(21) & \RegFile[7][22]~q\) ) ) ) # ( \RegFile[5][22]~q\ & ( !\R.curInst\(20) & ( 
-- (!\R.curInst\(21) & (\RegFile[4][22]~q\)) # (\R.curInst\(21) & ((\RegFile[6][22]~q\))) ) ) ) # ( !\RegFile[5][22]~q\ & ( !\R.curInst\(20) & ( (!\R.curInst\(21) & (\RegFile[4][22]~q\)) # (\R.curInst\(21) & ((\RegFile[6][22]~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100011101000111010001110100011100000000001100111100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[4][22]~q\,
	datab => \ALT_INV_R.curInst\(21),
	datac => \ALT_INV_RegFile[6][22]~q\,
	datad => \ALT_INV_RegFile[7][22]~q\,
	datae => \ALT_INV_RegFile[5][22]~q\,
	dataf => \ALT_INV_R.curInst\(20),
	combout => \Mux100~0_combout\);

-- Location: LABCELL_X62_Y1_N48
\Mux100~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux100~26_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (\R.curInst\(20) & (\RegFile[1][22]~q\))) # (\R.curInst\(22) & (((\Mux100~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (((\RegFile[2][22]~q\)))) # 
-- (\R.curInst\(20) & (\RegFile[3][22]~q\)))) # (\R.curInst\(22) & ((((\Mux100~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000000000111010000000000000011111111110001110111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[3][22]~q\,
	datab => \ALT_INV_R.curInst\(20),
	datac => \ALT_INV_RegFile[2][22]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux100~0_combout\,
	datag => \ALT_INV_RegFile[1][22]~q\,
	combout => \Mux100~26_combout\);

-- Location: LABCELL_X63_Y2_N6
\Mux100~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux100~13_combout\ = ( \Mux100~5_combout\ & ( \Mux100~26_combout\ & ( (!\R.curInst\(23)) # ((!\R.curInst\(24) & ((\Mux100~1_combout\))) # (\R.curInst\(24) & (\Mux100~9_combout\))) ) ) ) # ( !\Mux100~5_combout\ & ( \Mux100~26_combout\ & ( 
-- (!\R.curInst\(24) & (((!\R.curInst\(23)) # (\Mux100~1_combout\)))) # (\R.curInst\(24) & (\Mux100~9_combout\ & ((\R.curInst\(23))))) ) ) ) # ( \Mux100~5_combout\ & ( !\Mux100~26_combout\ & ( (!\R.curInst\(24) & (((\Mux100~1_combout\ & \R.curInst\(23))))) # 
-- (\R.curInst\(24) & (((!\R.curInst\(23))) # (\Mux100~9_combout\))) ) ) ) # ( !\Mux100~5_combout\ & ( !\Mux100~26_combout\ & ( (\R.curInst\(23) & ((!\R.curInst\(24) & ((\Mux100~1_combout\))) # (\R.curInst\(24) & (\Mux100~9_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110101000011110011010111110000001101011111111100110101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux100~9_combout\,
	datab => \ALT_INV_Mux100~1_combout\,
	datac => \ALT_INV_R.curInst\(24),
	datad => \ALT_INV_R.curInst\(23),
	datae => \ALT_INV_Mux100~5_combout\,
	dataf => \ALT_INV_Mux100~26_combout\,
	combout => \Mux100~13_combout\);

-- Location: MLABCELL_X72_Y4_N36
\NxR.aluData2[22]~28\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[22]~28_combout\ = ( \Equal4~1_combout\ & ( \Mux100~13_combout\ & ( (!\vAluSrc2~1_combout\) # (\Mux132~0_combout\) ) ) ) # ( !\Equal4~1_combout\ & ( \Mux100~13_combout\ & ( !\vAluSrc2~1_combout\ ) ) ) # ( \Equal4~1_combout\ & ( 
-- !\Mux100~13_combout\ & ( (\vAluSrc2~1_combout\ & \Mux132~0_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000110000001111001100110011001100111111001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_vAluSrc2~1_combout\,
	datac => \ALT_INV_Mux132~0_combout\,
	datae => \ALT_INV_Equal4~1_combout\,
	dataf => \ALT_INV_Mux100~13_combout\,
	combout => \NxR.aluData2[22]~28_combout\);

-- Location: FF_X72_Y4_N37
\R.aluData2[22]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR.aluData2[22]~28_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData2\(22));

-- Location: LABCELL_X77_Y7_N42
\ShiftRight0~12\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight0~12_combout\ = ( \ShiftRight1~31_OTERM45\ & ( (!\R.aluData2\(3) & (((!\R.aluData2\(2))) # (\ShiftRight1~32_OTERM21\))) # (\R.aluData2\(3) & (((\ShiftRight0~4_OTERM31\ & !\R.aluData2\(2))))) ) ) # ( !\ShiftRight1~31_OTERM45\ & ( 
-- (!\R.aluData2\(3) & (\ShiftRight1~32_OTERM21\ & ((\R.aluData2\(2))))) # (\R.aluData2\(3) & (((\ShiftRight0~4_OTERM31\ & !\R.aluData2\(2))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100100010000001010010001010101111001000101010111100100010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(3),
	datab => \ALT_INV_ShiftRight1~32_OTERM21\,
	datac => \ALT_INV_ShiftRight0~4_OTERM31\,
	datad => \ALT_INV_R.aluData2\(2),
	dataf => \ALT_INV_ShiftRight1~31_OTERM45\,
	combout => \ShiftRight0~12_combout\);

-- Location: LABCELL_X79_Y7_N24
\ShiftLeft0~39\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftLeft0~39_combout\ = ( \ShiftLeft0~22_OTERM737\ & ( \R.aluData2\(2) & ( (!\R.aluData2\(3) & ((\ShiftLeft0~30_OTERM601\))) # (\R.aluData2\(3) & (\ShiftLeft0~14_OTERM753\)) ) ) ) # ( !\ShiftLeft0~22_OTERM737\ & ( \R.aluData2\(2) & ( (!\R.aluData2\(3) & 
-- ((\ShiftLeft0~30_OTERM601\))) # (\R.aluData2\(3) & (\ShiftLeft0~14_OTERM753\)) ) ) ) # ( \ShiftLeft0~22_OTERM737\ & ( !\R.aluData2\(2) & ( (\R.aluData2\(3)) # (\ShiftLeft0~38_OTERM789\) ) ) ) # ( !\ShiftLeft0~22_OTERM737\ & ( !\R.aluData2\(2) & ( 
-- (\ShiftLeft0~38_OTERM789\ & !\R.aluData2\(3)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010100000000010101011111111100001111001100110000111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftLeft0~38_OTERM789\,
	datab => \ALT_INV_ShiftLeft0~14_OTERM753\,
	datac => \ALT_INV_ShiftLeft0~30_OTERM601\,
	datad => \ALT_INV_R.aluData2\(3),
	datae => \ALT_INV_ShiftLeft0~22_OTERM737\,
	dataf => \ALT_INV_R.aluData2\(2),
	combout => \ShiftLeft0~39_combout\);

-- Location: LABCELL_X80_Y9_N0
\Selector9~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector9~0_combout\ = ( \R.aluData2\(3) & ( \R.aluData1\(31) & ( \R.aluOp.ALUOpSRA~q\ ) ) ) # ( !\R.aluData2\(3) & ( \R.aluData1\(31) & ( (\R.aluOp.ALUOpSRA~q\ & ((!\R.aluData2\(2) & (\ShiftRight1~31_OTERM45\)) # (\R.aluData2\(2) & 
-- ((\ShiftRight1~32_OTERM21\))))) ) ) ) # ( !\R.aluData2\(3) & ( !\R.aluData1\(31) & ( (\R.aluOp.ALUOpSRA~q\ & ((!\R.aluData2\(2) & (\ShiftRight1~31_OTERM45\)) # (\R.aluData2\(2) & ((\ShiftRight1~32_OTERM21\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010000000111000000000000000000000100000001110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~31_OTERM45\,
	datab => \ALT_INV_R.aluData2\(2),
	datac => \ALT_INV_R.aluOp.ALUOpSRA~q\,
	datad => \ALT_INV_ShiftRight1~32_OTERM21\,
	datae => \ALT_INV_R.aluData2\(3),
	dataf => \ALT_INV_R.aluData1\(31),
	combout => \Selector9~0_combout\);

-- Location: LABCELL_X81_Y7_N24
\Selector9~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector9~1_combout\ = ( !\R.aluData2\(4) & ( \Selector9~0_combout\ ) ) # ( !\R.aluData2\(4) & ( !\Selector9~0_combout\ & ( (!\ShiftRight0~12_combout\ & (\ShiftLeft0~39_combout\ & ((\R.aluOp.ALUOpSLL~q\)))) # (\ShiftRight0~12_combout\ & 
-- (((\ShiftLeft0~39_combout\ & \R.aluOp.ALUOpSLL~q\)) # (\R.aluOp.ALUOpSRL~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100110111000000000000000011111111111111110000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight0~12_combout\,
	datab => \ALT_INV_ShiftLeft0~39_combout\,
	datac => \ALT_INV_R.aluOp.ALUOpSRL~q\,
	datad => \ALT_INV_R.aluOp.ALUOpSLL~q\,
	datae => \ALT_INV_R.aluData2\(4),
	dataf => \ALT_INV_Selector9~0_combout\,
	combout => \Selector9~1_combout\);

-- Location: LABCELL_X77_Y8_N9
\Selector9~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector9~3_combout\ = ( \R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( (!\R.aluOp.ALUOpOr~q\ & (\R.aluData2\(23) & \R.aluData1\(23))) # (\R.aluOp.ALUOpOr~q\ & ((\R.aluData1\(23)) # (\R.aluData2\(23)))) ) ) # ( !\R.aluOp.ALUOpAnd~DUPLICATE_q\ & ( 
-- (\R.aluOp.ALUOpOr~q\ & ((\R.aluData1\(23)) # (\R.aluData2\(23)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100110011000000110011001100000011001111110000001100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluOp.ALUOpOr~q\,
	datac => \ALT_INV_R.aluData2\(23),
	datad => \ALT_INV_R.aluData1\(23),
	dataf => \ALT_INV_R.aluOp.ALUOpAnd~DUPLICATE_q\,
	combout => \Selector9~3_combout\);

-- Location: LABCELL_X75_Y5_N12
\LessThan1~30\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~30_combout\ = ( \Mux131~0_combout\ & ( \Mux99~13_combout\ & ( !\Mux231~0_combout\ $ (((!\Equal4~1_combout\ & \vAluSrc2~1_combout\))) ) ) ) # ( !\Mux131~0_combout\ & ( \Mux99~13_combout\ & ( !\vAluSrc2~1_combout\ $ (\Mux231~0_combout\) ) ) ) # ( 
-- \Mux131~0_combout\ & ( !\Mux99~13_combout\ & ( !\Mux231~0_combout\ $ (((!\Equal4~1_combout\) # (!\vAluSrc2~1_combout\))) ) ) ) # ( !\Mux131~0_combout\ & ( !\Mux99~13_combout\ & ( \Mux231~0_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111000100011110111011001100001100111101110100100010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Equal4~1_combout\,
	datab => \ALT_INV_vAluSrc2~1_combout\,
	datad => \ALT_INV_Mux231~0_combout\,
	datae => \ALT_INV_Mux131~0_combout\,
	dataf => \ALT_INV_Mux99~13_combout\,
	combout => \LessThan1~30_combout\);

-- Location: FF_X75_Y5_N13
\LessThan1~30_NEW_REG42\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \LessThan1~30_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \LessThan1~30_OTERM43\);

-- Location: LABCELL_X77_Y8_N12
\Selector9~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector9~2_combout\ = ( \ShiftLeft0~9_OTERM461\ & ( (\Selector12~2_OTERM395\ & (!\R.aluData2\(3) & ((!\R.aluData2\(2)) # (\ShiftLeft0~3_OTERM223\)))) ) ) # ( !\ShiftLeft0~9_OTERM461\ & ( (\Selector12~2_OTERM395\ & (\ShiftLeft0~3_OTERM223\ & 
-- (!\R.aluData2\(3) & \R.aluData2\(2)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000010000000000000001000001010000000100000101000000010000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector12~2_OTERM395\,
	datab => \ALT_INV_ShiftLeft0~3_OTERM223\,
	datac => \ALT_INV_R.aluData2\(3),
	datad => \ALT_INV_R.aluData2\(2),
	dataf => \ALT_INV_ShiftLeft0~9_OTERM461\,
	combout => \Selector9~2_combout\);

-- Location: LABCELL_X77_Y8_N0
\Selector9~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector9~4_combout\ = ( !\Selector9~2_combout\ & ( (!\Selector17~0_OTERM391\ & (!\Selector9~3_combout\ & ((!\LessThan1~30_OTERM43\) # (!\R.aluOp.ALUOpXor~DUPLICATE_q\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000100010000000100010001000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector17~0_OTERM391\,
	datab => \ALT_INV_Selector9~3_combout\,
	datac => \ALT_INV_LessThan1~30_OTERM43\,
	datad => \ALT_INV_R.aluOp.ALUOpXor~DUPLICATE_q\,
	dataf => \ALT_INV_Selector9~2_combout\,
	combout => \Selector9~4_combout\);

-- Location: LABCELL_X80_Y4_N6
\Selector9~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector9~5_combout\ = ( \Add2~93_sumout\ & ( \Selector9~4_combout\ & ( (((\R.aluOp.ALUOpAdd~q\ & \Add1~93_sumout\)) # (\Selector9~1_combout\)) # (\R.aluOp.ALUOpSub~q\) ) ) ) # ( !\Add2~93_sumout\ & ( \Selector9~4_combout\ & ( ((\R.aluOp.ALUOpAdd~q\ & 
-- \Add1~93_sumout\)) # (\Selector9~1_combout\) ) ) ) # ( \Add2~93_sumout\ & ( !\Selector9~4_combout\ ) ) # ( !\Add2~93_sumout\ & ( !\Selector9~4_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111111111111111111100000011111111110101011111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datab => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datac => \ALT_INV_Add1~93_sumout\,
	datad => \ALT_INV_Selector9~1_combout\,
	datae => \ALT_INV_Add2~93_sumout\,
	dataf => \ALT_INV_Selector9~4_combout\,
	combout => \Selector9~5_combout\);

-- Location: LABCELL_X80_Y4_N0
\Comb:vJumpAdr[23]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[23]~0_combout\ = ( \R.aluRes\(23) & ( \Add3~93_sumout\ & ( ((!\R.aluCalc~q\) # (!\Equal4~2_combout\)) # (\Selector9~5_combout\) ) ) ) # ( !\R.aluRes\(23) & ( \Add3~93_sumout\ & ( (!\Equal4~2_combout\) # ((\Selector9~5_combout\ & 
-- \R.aluCalc~q\)) ) ) ) # ( \R.aluRes\(23) & ( !\Add3~93_sumout\ & ( (\Equal4~2_combout\ & ((!\R.aluCalc~q\) # (\Selector9~5_combout\))) ) ) ) # ( !\R.aluRes\(23) & ( !\Add3~93_sumout\ & ( (\Selector9~5_combout\ & (\R.aluCalc~q\ & \Equal4~2_combout\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000011000000001111001111111111000000111111111111110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Selector9~5_combout\,
	datac => \ALT_INV_R.aluCalc~q\,
	datad => \ALT_INV_Equal4~2_combout\,
	datae => \ALT_INV_R.aluRes\(23),
	dataf => \ALT_INV_Add3~93_sumout\,
	combout => \Comb:vJumpAdr[23]~0_combout\);

-- Location: FF_X80_Y4_N1
\R.curPC[23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[23]~0_combout\,
	asdata => \Add0~85_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(23));

-- Location: IOIBUF_X36_Y0_N1
\avm_d_readdata[15]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_readdata(15),
	o => \avm_d_readdata[15]~input_o\);

-- Location: MLABCELL_X78_Y5_N54
\Comb:vRegWriteData[23]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[23]~1_combout\ = ( \R.curInst\(13) & ( \Add1~93_sumout\ & ( (!\R.memToReg~q\ & (((\R.aluOp.ALUOpAdd~q\)))) # (\R.memToReg~q\ & (!\R.curInst\(14) & ((\avm_d_readdata[15]~input_o\)))) ) ) ) # ( !\R.curInst\(13) & ( \Add1~93_sumout\ & ( 
-- (!\R.memToReg~q\ & ((\R.aluOp.ALUOpAdd~q\))) # (\R.memToReg~q\ & (!\R.curInst\(14))) ) ) ) # ( \R.curInst\(13) & ( !\Add1~93_sumout\ & ( (!\R.curInst\(14) & (\R.memToReg~q\ & \avm_d_readdata[15]~input_o\)) ) ) ) # ( !\R.curInst\(13) & ( !\Add1~93_sumout\ 
-- & ( (!\R.curInst\(14) & \R.memToReg~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101000001010000000000000101000111010001110100011000000111010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(14),
	datab => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datac => \ALT_INV_R.memToReg~q\,
	datad => \ALT_INV_avm_d_readdata[15]~input_o\,
	datae => \ALT_INV_R.curInst\(13),
	dataf => \ALT_INV_Add1~93_sumout\,
	combout => \Comb:vRegWriteData[23]~1_combout\);

-- Location: LABCELL_X80_Y4_N27
\Comb:vRegWriteData[23]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[23]~3_combout\ = ( \Selector9~4_combout\ & ( (!\R.aluCalc~q\ & (!\R.memToReg~q\ & ((!\R.aluRes\(23))))) # (\R.aluCalc~q\ & (((!\Selector9~1_combout\)))) ) ) # ( !\Selector9~4_combout\ & ( (!\R.memToReg~q\ & (!\R.aluCalc~q\ & 
-- !\R.aluRes\(23))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000100000000000100010000000000010111000001100001011100000110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.memToReg~q\,
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_Selector9~1_combout\,
	datad => \ALT_INV_R.aluRes\(23),
	dataf => \ALT_INV_Selector9~4_combout\,
	combout => \Comb:vRegWriteData[23]~3_combout\);

-- Location: LABCELL_X79_Y1_N18
\Comb:vRegWriteData[23]~2_RESYN1114\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[23]~2_RESYN1114_BDD1115\ = ( \R.curInst\(12) & ( !\avm_d_readdata[23]~input_o\ ) ) # ( !\R.curInst\(12) & ( !\avm_d_readdata[31]~input_o\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010101010101010101010101010101011110000111100001111000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_avm_d_readdata[31]~input_o\,
	datac => \ALT_INV_avm_d_readdata[23]~input_o\,
	dataf => \ALT_INV_R.curInst\(12),
	combout => \Comb:vRegWriteData[23]~2_RESYN1114_BDD1115\);

-- Location: LABCELL_X79_Y1_N39
\Comb:vRegWriteData[23]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[23]~2_combout\ = ( \R.curInst\(13) & ( \Comb:vRegWriteData[23]~2_RESYN1114_BDD1115\ & ( (\R.memToReg~q\ & (((!\avm_d_readdata[15]~input_o\) # (\R.curInst\(14))) # (\R.curInst\(12)))) ) ) ) # ( !\R.curInst\(13) & ( 
-- \Comb:vRegWriteData[23]~2_RESYN1114_BDD1115\ & ( \R.memToReg~q\ ) ) ) # ( \R.curInst\(13) & ( !\Comb:vRegWriteData[23]~2_RESYN1114_BDD1115\ & ( (\R.memToReg~q\ & (((!\avm_d_readdata[15]~input_o\) # (\R.curInst\(14))) # (\R.curInst\(12)))) ) ) ) # ( 
-- !\R.curInst\(13) & ( !\Comb:vRegWriteData[23]~2_RESYN1114_BDD1115\ & ( (\R.memToReg~q\ & \R.curInst\(14)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000001111000011010000111100001111000011110000110100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(12),
	datab => \ALT_INV_avm_d_readdata[15]~input_o\,
	datac => \ALT_INV_R.memToReg~q\,
	datad => \ALT_INV_R.curInst\(14),
	datae => \ALT_INV_R.curInst\(13),
	dataf => \ALT_INV_Comb:vRegWriteData[23]~2_RESYN1114_BDD1115\,
	combout => \Comb:vRegWriteData[23]~2_combout\);

-- Location: LABCELL_X81_Y5_N0
\Comb:vRegWriteData[23]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[23]~0_combout\ = ( !\Comb:vRegWriteData[23]~2_combout\ & ( \Add2~93_sumout\ & ( (!\Comb:vRegWriteData[23]~3_combout\) # ((\R.aluCalc~q\ & ((\R.aluOp.ALUOpSub~q\) # (\Comb:vRegWriteData[23]~1_combout\)))) ) ) ) # ( 
-- !\Comb:vRegWriteData[23]~2_combout\ & ( !\Add2~93_sumout\ & ( (!\Comb:vRegWriteData[23]~3_combout\) # ((\Comb:vRegWriteData[23]~1_combout\ & \R.aluCalc~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111000011110101000000000000000011110000111101110000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Comb:vRegWriteData[23]~1_combout\,
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datac => \ALT_INV_Comb:vRegWriteData[23]~3_combout\,
	datad => \ALT_INV_R.aluCalc~q\,
	datae => \ALT_INV_Comb:vRegWriteData[23]~2_combout\,
	dataf => \ALT_INV_Add2~93_sumout\,
	combout => \Comb:vRegWriteData[23]~0_combout\);

-- Location: FF_X81_Y5_N35
\R.regWriteData[23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Add0~85_sumout\,
	asdata => \Comb:vRegWriteData[23]~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(23));

-- Location: FF_X68_Y2_N56
\RegFile[15][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(23),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~8_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[15][23]~q\);

-- Location: LABCELL_X68_Y2_N30
\Mux99~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux99~14_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & (\RegFile[8][23]~q\)) # (\R.curInst\(20) & ((\RegFile[9][23]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & ((\RegFile[10][23]~q\))) # (\R.curInst\(20) & (\RegFile[11][23]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110000110011111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[11][23]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[10][23]~q\,
	datad => \ALT_INV_RegFile[9][23]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][23]~q\,
	combout => \Mux99~14_combout\);

-- Location: LABCELL_X62_Y2_N30
\Mux99~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux99~1_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux99~14_combout\)))) # (\R.curInst\(22) & ((!\Mux99~14_combout\ & (\RegFile[12][23]~q\)) # (\Mux99~14_combout\ & ((\RegFile[13][23]~q\)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) 
-- & ((((\Mux99~14_combout\))))) # (\R.curInst\(22) & (((!\Mux99~14_combout\ & ((\RegFile[14][23]~q\))) # (\Mux99~14_combout\ & (\RegFile[15][23]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111001100111111111101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][23]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[14][23]~q\,
	datad => \ALT_INV_RegFile[13][23]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux99~14_combout\,
	datag => \ALT_INV_RegFile[12][23]~q\,
	combout => \Mux99~1_combout\);

-- Location: FF_X64_Y1_N23
\RegFile[16][23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[16][23]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~25_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[16][23]~q\);

-- Location: LABCELL_X64_Y1_N24
\Mux99~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux99~18_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[16][23]~q\))) # (\R.curInst\(20) & (\RegFile[17][23]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & (\RegFile[18][23]~q\)) # (\R.curInst\(20) & ((\RegFile[19][23]~q\)))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001110111011101110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[17][23]~q\,
	datac => \ALT_INV_RegFile[18][23]~q\,
	datad => \ALT_INV_RegFile[19][23]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][23]~q\,
	combout => \Mux99~18_combout\);

-- Location: LABCELL_X64_Y1_N48
\Mux99~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux99~5_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux99~18_combout\)))) # (\R.curInst\(22) & ((!\Mux99~18_combout\ & ((\RegFile[20][23]~q\))) # (\Mux99~18_combout\ & (\RegFile[21][23]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux99~18_combout\)))) # (\R.curInst\(22) & ((!\Mux99~18_combout\ & ((\RegFile[22][23]~q\))) # (\Mux99~18_combout\ & (\RegFile[23][23]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111010101011111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][23]~q\,
	datab => \ALT_INV_RegFile[23][23]~q\,
	datac => \ALT_INV_RegFile[22][23]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux99~18_combout\,
	datag => \ALT_INV_RegFile[20][23]~q\,
	combout => \Mux99~5_combout\);

-- Location: LABCELL_X63_Y2_N12
\Mux99~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux99~22_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & (\RegFile[24][23]~q\)) # (\R.curInst\(20) & ((\RegFile[25][23]~q\)))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & ((\RegFile[26][23]~q\))) # (\R.curInst\(20) & (\RegFile[27][23]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000101000001010000010100000101001010101111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[27][23]~q\,
	datac => \ALT_INV_RegFile[26][23]~q\,
	datad => \ALT_INV_RegFile[25][23]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][23]~q\,
	combout => \Mux99~22_combout\);

-- Location: LABCELL_X63_Y2_N54
\Mux99~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux99~9_combout\ = ( !\R.curInst\(21) & ( ((!\Mux99~22_combout\ & (\RegFile[28][23]~q\ & ((\R.curInst\(22))))) # (\Mux99~22_combout\ & (((!\R.curInst\(22)) # (\RegFile[29][23]~q\))))) ) ) # ( \R.curInst\(21) & ( (!\Mux99~22_combout\ & 
-- (((\RegFile[30][23]~q\ & ((\R.curInst\(22))))))) # (\Mux99~22_combout\ & ((((!\R.curInst\(22)))) # (\RegFile[31][23]~q\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0011001100110011001100110011001100001100001111110001110100011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[31][23]~q\,
	datab => \ALT_INV_Mux99~22_combout\,
	datac => \ALT_INV_RegFile[30][23]~q\,
	datad => \ALT_INV_RegFile[29][23]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(22),
	datag => \ALT_INV_RegFile[28][23]~q\,
	combout => \Mux99~9_combout\);

-- Location: LABCELL_X73_Y3_N24
\Mux99~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux99~0_combout\ = ( \RegFile[6][23]~q\ & ( \R.curInst\(20) & ( (!\R.curInst\(21) & (\RegFile[5][23]~q\)) # (\R.curInst\(21) & ((\RegFile[7][23]~q\))) ) ) ) # ( !\RegFile[6][23]~q\ & ( \R.curInst\(20) & ( (!\R.curInst\(21) & (\RegFile[5][23]~q\)) # 
-- (\R.curInst\(21) & ((\RegFile[7][23]~q\))) ) ) ) # ( \RegFile[6][23]~q\ & ( !\R.curInst\(20) & ( (\R.curInst\(21)) # (\RegFile[4][23]~q\) ) ) ) # ( !\RegFile[6][23]~q\ & ( !\R.curInst\(20) & ( (\RegFile[4][23]~q\ & !\R.curInst\(21)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011000000110000001111110011111101010000010111110101000001011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[5][23]~q\,
	datab => \ALT_INV_RegFile[4][23]~q\,
	datac => \ALT_INV_R.curInst\(21),
	datad => \ALT_INV_RegFile[7][23]~q\,
	datae => \ALT_INV_RegFile[6][23]~q\,
	dataf => \ALT_INV_R.curInst\(20),
	combout => \Mux99~0_combout\);

-- Location: LABCELL_X62_Y1_N6
\Mux99~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux99~26_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (\R.curInst\(20) & (\RegFile[1][23]~q\))) # (\R.curInst\(22) & (((\Mux99~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (((\RegFile[2][23]~q\)))) # 
-- (\R.curInst\(20) & (\RegFile[3][23]~q\)))) # (\R.curInst\(22) & ((((\Mux99~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000010100000000000110110000000000000101111111110001101111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(20),
	datab => \ALT_INV_RegFile[3][23]~q\,
	datac => \ALT_INV_RegFile[2][23]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux99~0_combout\,
	datag => \ALT_INV_RegFile[1][23]~q\,
	combout => \Mux99~26_combout\);

-- Location: LABCELL_X63_Y2_N48
\Mux99~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux99~13_combout\ = ( \Mux99~9_combout\ & ( \Mux99~26_combout\ & ( (!\R.curInst\(24) & ((!\R.curInst\(23)) # ((\Mux99~1_combout\)))) # (\R.curInst\(24) & (((\Mux99~5_combout\)) # (\R.curInst\(23)))) ) ) ) # ( !\Mux99~9_combout\ & ( \Mux99~26_combout\ & ( 
-- (!\R.curInst\(24) & ((!\R.curInst\(23)) # ((\Mux99~1_combout\)))) # (\R.curInst\(24) & (!\R.curInst\(23) & ((\Mux99~5_combout\)))) ) ) ) # ( \Mux99~9_combout\ & ( !\Mux99~26_combout\ & ( (!\R.curInst\(24) & (\R.curInst\(23) & (\Mux99~1_combout\))) # 
-- (\R.curInst\(24) & (((\Mux99~5_combout\)) # (\R.curInst\(23)))) ) ) ) # ( !\Mux99~9_combout\ & ( !\Mux99~26_combout\ & ( (!\R.curInst\(24) & (\R.curInst\(23) & (\Mux99~1_combout\))) # (\R.curInst\(24) & (!\R.curInst\(23) & ((\Mux99~5_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001001000110000100110101011110001010110011101001101111011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(24),
	datab => \ALT_INV_R.curInst\(23),
	datac => \ALT_INV_Mux99~1_combout\,
	datad => \ALT_INV_Mux99~5_combout\,
	datae => \ALT_INV_Mux99~9_combout\,
	dataf => \ALT_INV_Mux99~26_combout\,
	combout => \Mux99~13_combout\);

-- Location: LABCELL_X75_Y5_N30
\NxR.aluData2[23]~27\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[23]~27_combout\ = ( \Mux131~0_combout\ & ( \Mux99~13_combout\ & ( (!\vAluSrc2~1_combout\) # (\Equal4~1_combout\) ) ) ) # ( !\Mux131~0_combout\ & ( \Mux99~13_combout\ & ( !\vAluSrc2~1_combout\ ) ) ) # ( \Mux131~0_combout\ & ( 
-- !\Mux99~13_combout\ & ( (\Equal4~1_combout\ & \vAluSrc2~1_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000100010001000111001100110011001101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Equal4~1_combout\,
	datab => \ALT_INV_vAluSrc2~1_combout\,
	datae => \ALT_INV_Mux131~0_combout\,
	dataf => \ALT_INV_Mux99~13_combout\,
	combout => \NxR.aluData2[23]~27_combout\);

-- Location: FF_X75_Y5_N31
\R.aluData2[23]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR.aluData2[23]~27_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData2\(23));

-- Location: LABCELL_X61_Y5_N30
\LessThan1~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~29_combout\ = ( \Mux130~0_combout\ & ( \Mux230~0_combout\ & ( (!\vAluSrc2~1_combout\ & (!\Mux98~13_combout\)) # (\vAluSrc2~1_combout\ & ((!\Equal4~1_combout\))) ) ) ) # ( !\Mux130~0_combout\ & ( \Mux230~0_combout\ & ( (!\Mux98~13_combout\) # 
-- (\vAluSrc2~1_combout\) ) ) ) # ( \Mux130~0_combout\ & ( !\Mux230~0_combout\ & ( (!\vAluSrc2~1_combout\ & (\Mux98~13_combout\)) # (\vAluSrc2~1_combout\ & ((\Equal4~1_combout\))) ) ) ) # ( !\Mux130~0_combout\ & ( !\Mux230~0_combout\ & ( (\Mux98~13_combout\ 
-- & !\vAluSrc2~1_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011000000110000001100000011111111001111110011111100111111000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Mux98~13_combout\,
	datac => \ALT_INV_vAluSrc2~1_combout\,
	datad => \ALT_INV_Equal4~1_combout\,
	datae => \ALT_INV_Mux130~0_combout\,
	dataf => \ALT_INV_Mux230~0_combout\,
	combout => \LessThan1~29_combout\);

-- Location: FF_X61_Y5_N31
\LessThan1~29_NEW_REG46\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \LessThan1~29_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \LessThan1~29_OTERM47\);

-- Location: FF_X79_Y5_N55
\R.aluData2[25]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR.aluData2[25]~22_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData2\(25));

-- Location: LABCELL_X73_Y4_N18
\LessThan1~28_RTM053\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~28_RTM053_combout\ = ( \Mux227~0_combout\ & ( \NxR.aluData2[28]~23_combout\ & ( (!\NxR.aluData2[27]~24_combout\) # ((!\Mux226~0_combout\) # (!\Mux228~0_combout\ $ (!\NxR.aluData2[26]~25_combout\))) ) ) ) # ( !\Mux227~0_combout\ & ( 
-- \NxR.aluData2[28]~23_combout\ & ( ((!\Mux226~0_combout\) # (!\Mux228~0_combout\ $ (!\NxR.aluData2[26]~25_combout\))) # (\NxR.aluData2[27]~24_combout\) ) ) ) # ( \Mux227~0_combout\ & ( !\NxR.aluData2[28]~23_combout\ & ( (!\NxR.aluData2[27]~24_combout\) # 
-- ((!\Mux228~0_combout\ $ (!\NxR.aluData2[26]~25_combout\)) # (\Mux226~0_combout\)) ) ) ) # ( !\Mux227~0_combout\ & ( !\NxR.aluData2[28]~23_combout\ & ( ((!\Mux228~0_combout\ $ (!\NxR.aluData2[26]~25_combout\)) # (\Mux226~0_combout\)) # 
-- (\NxR.aluData2[27]~24_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0111110111111111101111101111111111111111011111011111111110111110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_NxR.aluData2[27]~24_combout\,
	datab => \ALT_INV_Mux228~0_combout\,
	datac => \ALT_INV_NxR.aluData2[26]~25_combout\,
	datad => \ALT_INV_Mux226~0_combout\,
	datae => \ALT_INV_Mux227~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[28]~23_combout\,
	combout => \LessThan1~28_RTM053_combout\);

-- Location: FF_X73_Y4_N19
\LessThan1~28_NEW_REG50\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \LessThan1~28_RTM053_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \LessThan1~28_OTERM51\);

-- Location: LABCELL_X80_Y5_N18
\LessThan1~33\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~33_combout\ = ( \R.aluData1\(25) & ( (!\LessThan1~29_OTERM47\ & (\R.aluData2\(25) & !\LessThan1~28_OTERM51\)) ) ) # ( !\R.aluData1\(25) & ( (!\LessThan1~29_OTERM47\ & (!\R.aluData2\(25) & !\LessThan1~28_OTERM51\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1100000000000000110000000000000000001100000000000000110000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_LessThan1~29_OTERM47\,
	datac => \ALT_INV_R.aluData2\(25),
	datad => \ALT_INV_LessThan1~28_OTERM51\,
	dataf => \ALT_INV_R.aluData1\(25),
	combout => \LessThan1~33_combout\);

-- Location: LABCELL_X73_Y4_N12
\LessThan1~34\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~34_combout\ = ( \NxR.aluData2[26]~25_combout\ & ( \Mux228~0_combout\ & ( (!\Mux226~0_combout\ & (((\NxR.aluData2[27]~24_combout\ & !\Mux227~0_combout\)) # (\NxR.aluData2[28]~23_combout\))) # (\Mux226~0_combout\ & (\NxR.aluData2[27]~24_combout\ 
-- & (\NxR.aluData2[28]~23_combout\ & !\Mux227~0_combout\))) ) ) ) # ( !\NxR.aluData2[26]~25_combout\ & ( \Mux228~0_combout\ & ( (!\Mux226~0_combout\ & (((\NxR.aluData2[27]~24_combout\ & !\Mux227~0_combout\)) # (\NxR.aluData2[28]~23_combout\))) # 
-- (\Mux226~0_combout\ & (\NxR.aluData2[27]~24_combout\ & (\NxR.aluData2[28]~23_combout\ & !\Mux227~0_combout\))) ) ) ) # ( \NxR.aluData2[26]~25_combout\ & ( !\Mux228~0_combout\ & ( (!\Mux226~0_combout\ & (((!\Mux227~0_combout\) # 
-- (\NxR.aluData2[28]~23_combout\)) # (\NxR.aluData2[27]~24_combout\))) # (\Mux226~0_combout\ & (\NxR.aluData2[28]~23_combout\ & ((!\Mux227~0_combout\) # (\NxR.aluData2[27]~24_combout\)))) ) ) ) # ( !\NxR.aluData2[26]~25_combout\ & ( !\Mux228~0_combout\ & ( 
-- (!\Mux226~0_combout\ & (((\NxR.aluData2[27]~24_combout\ & !\Mux227~0_combout\)) # (\NxR.aluData2[28]~23_combout\))) # (\Mux226~0_combout\ & (\NxR.aluData2[27]~24_combout\ & (\NxR.aluData2[28]~23_combout\ & !\Mux227~0_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100110100001100110011110100110101001101000011000100110100001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_NxR.aluData2[27]~24_combout\,
	datab => \ALT_INV_Mux226~0_combout\,
	datac => \ALT_INV_NxR.aluData2[28]~23_combout\,
	datad => \ALT_INV_Mux227~0_combout\,
	datae => \ALT_INV_NxR.aluData2[26]~25_combout\,
	dataf => \ALT_INV_Mux228~0_combout\,
	combout => \LessThan1~34_combout\);

-- Location: FF_X73_Y4_N13
\LessThan1~34_NEW_REG54\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \LessThan1~34_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \LessThan1~34_OTERM55\);

-- Location: MLABCELL_X84_Y5_N36
\LessThan1~35\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~35_combout\ = ( \R.aluData1\(25) & ( !\LessThan1~34_OTERM55\ & ( ((!\R.aluData2\(24)) # ((!\R.aluData2\(25)) # (\LessThan1~28_OTERM51\))) # (\R.aluData1\(24)) ) ) ) # ( !\R.aluData1\(25) & ( !\LessThan1~34_OTERM55\ & ( ((!\R.aluData2\(25) & 
-- ((!\R.aluData2\(24)) # (\R.aluData1\(24))))) # (\LessThan1~28_OTERM51\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1101000011111111111111011111111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData1\(24),
	datab => \ALT_INV_R.aluData2\(24),
	datac => \ALT_INV_R.aluData2\(25),
	datad => \ALT_INV_LessThan1~28_OTERM51\,
	datae => \ALT_INV_R.aluData1\(25),
	dataf => \ALT_INV_LessThan1~34_OTERM55\,
	combout => \LessThan1~35_combout\);

-- Location: LABCELL_X80_Y5_N36
\LessThan1~36\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~36_combout\ = ( \R.aluData2\(22) & ( \R.aluData1\(22) & ( (\LessThan1~35_combout\ & ((!\R.aluData2\(23)) # ((!\LessThan1~33_combout\) # (\R.aluData1\(23))))) ) ) ) # ( !\R.aluData2\(22) & ( \R.aluData1\(22) & ( (\LessThan1~35_combout\ & 
-- ((!\R.aluData2\(23)) # ((!\LessThan1~33_combout\) # (\R.aluData1\(23))))) ) ) ) # ( \R.aluData2\(22) & ( !\R.aluData1\(22) & ( (\LessThan1~35_combout\ & ((!\LessThan1~33_combout\) # ((!\R.aluData2\(23) & \R.aluData1\(23))))) ) ) ) # ( !\R.aluData2\(22) & 
-- ( !\R.aluData1\(22) & ( (\LessThan1~35_combout\ & ((!\R.aluData2\(23)) # ((!\LessThan1~33_combout\) # (\R.aluData1\(23))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111011000000001111001000000000111110110000000011111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(23),
	datab => \ALT_INV_R.aluData1\(23),
	datac => \ALT_INV_LessThan1~33_combout\,
	datad => \ALT_INV_LessThan1~35_combout\,
	datae => \ALT_INV_R.aluData2\(22),
	dataf => \ALT_INV_R.aluData1\(22),
	combout => \LessThan1~36_combout\);

-- Location: LABCELL_X81_Y7_N6
\LessThan1~38\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~38_combout\ = ( \R.aluData2\(31) & ( \R.aluData2\(30) & ( (\R.aluData1\(31) & ((!\R.aluData1\(30)) # ((!\R.aluData1\(29) & \R.aluData2\(29))))) ) ) ) # ( !\R.aluData2\(31) & ( \R.aluData2\(30) & ( (!\R.aluData1\(31) & ((!\R.aluData1\(30)) # 
-- ((!\R.aluData1\(29) & \R.aluData2\(29))))) ) ) ) # ( \R.aluData2\(31) & ( !\R.aluData2\(30) & ( (!\R.aluData1\(30) & (!\R.aluData1\(29) & (\R.aluData2\(29) & \R.aluData1\(31)))) ) ) ) # ( !\R.aluData2\(31) & ( !\R.aluData2\(30) & ( (!\R.aluData1\(30) & 
-- (!\R.aluData1\(29) & (\R.aluData2\(29) & !\R.aluData1\(31)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000100000000000000000000000100010101110000000000000000010101110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData1\(30),
	datab => \ALT_INV_R.aluData1\(29),
	datac => \ALT_INV_R.aluData2\(29),
	datad => \ALT_INV_R.aluData1\(31),
	datae => \ALT_INV_R.aluData2\(31),
	dataf => \ALT_INV_R.aluData2\(30),
	combout => \LessThan1~38_combout\);

-- Location: LABCELL_X81_Y7_N48
\LessThan1~37\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~37_combout\ = ( \R.aluData1\(30) & ( \R.aluData2\(30) & ( (!\R.aluData2\(31) & (!\R.aluData1\(31) & (!\R.aluData1\(29) $ (\R.aluData2\(29))))) # (\R.aluData2\(31) & (\R.aluData1\(31) & (!\R.aluData1\(29) $ (\R.aluData2\(29))))) ) ) ) # ( 
-- !\R.aluData1\(30) & ( !\R.aluData2\(30) & ( (!\R.aluData2\(31) & (!\R.aluData1\(31) & (!\R.aluData1\(29) $ (\R.aluData2\(29))))) # (\R.aluData2\(31) & (\R.aluData1\(31) & (!\R.aluData1\(29) $ (\R.aluData2\(29))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000001001000001000000000000000000000000000000001000001001000001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(31),
	datab => \ALT_INV_R.aluData1\(29),
	datac => \ALT_INV_R.aluData2\(29),
	datad => \ALT_INV_R.aluData1\(31),
	datae => \ALT_INV_R.aluData1\(30),
	dataf => \ALT_INV_R.aluData2\(30),
	combout => \LessThan1~37_combout\);

-- Location: LABCELL_X75_Y5_N54
\Mux20~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux20~0_combout\ = ( \R.curInst\(14) & ( \R.curInst\(13) & ( (\R.aluOp.ALUOpSLTU~q\ & \R.curInst\(6)) ) ) ) # ( !\R.curInst\(14) & ( \R.curInst\(13) & ( (!\R.curInst\(6) & (\R.curInst\(12) & ((!\R.curInst\(2))))) # (\R.curInst\(6) & 
-- (((\R.aluOp.ALUOpSLTU~q\)))) ) ) ) # ( \R.curInst\(14) & ( !\R.curInst\(13) & ( (\R.aluOp.ALUOpSLTU~q\ & \R.curInst\(6)) ) ) ) # ( !\R.curInst\(14) & ( !\R.curInst\(13) & ( (\R.aluOp.ALUOpSLTU~q\ & \R.curInst\(6)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110011000000000011001101010000001100110000000000110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(12),
	datab => \ALT_INV_R.aluOp.ALUOpSLTU~q\,
	datac => \ALT_INV_R.curInst\(2),
	datad => \ALT_INV_R.curInst\(6),
	datae => \ALT_INV_R.curInst\(14),
	dataf => \ALT_INV_R.curInst\(13),
	combout => \Mux20~0_combout\);

-- Location: LABCELL_X77_Y6_N57
\Mux20~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux20~1_combout\ = ( \R.aluOp.ALUOpSLTU~q\ & ( \Mux20~0_combout\ & ( ((!\R.curInst\(3) & (!\Mux26~0_combout\)) # (\R.curInst\(3) & ((!\Mux123~0_combout\)))) # (\R.curInst\(4)) ) ) ) # ( !\R.aluOp.ALUOpSLTU~q\ & ( \Mux20~0_combout\ & ( (!\R.curInst\(3) & 
-- \R.curInst\(4)) ) ) ) # ( \R.aluOp.ALUOpSLTU~q\ & ( !\Mux20~0_combout\ & ( (!\R.curInst\(3) & (!\Mux26~0_combout\ & ((!\R.curInst\(4))))) # (\R.curInst\(3) & (((!\Mux123~0_combout\) # (\R.curInst\(4))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110110000101010100000000101010101101100011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(3),
	datab => \ALT_INV_Mux26~0_combout\,
	datac => \ALT_INV_Mux123~0_combout\,
	datad => \ALT_INV_R.curInst\(4),
	datae => \ALT_INV_R.aluOp.ALUOpSLTU~q\,
	dataf => \ALT_INV_Mux20~0_combout\,
	combout => \Mux20~1_combout\);

-- Location: LABCELL_X75_Y5_N42
\R.aluOp.ALUOpSLTU_NEW570\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.aluOp.ALUOpSLTU_OTERM571\ = ( \R.aluOp.ALUOpSLTU~q\ & ( \Mux20~1_combout\ ) ) # ( !\R.aluOp.ALUOpSLTU~q\ & ( \Mux20~1_combout\ & ( \vAluSrc2~0_combout\ ) ) ) # ( \R.aluOp.ALUOpSLTU~q\ & ( !\Mux20~1_combout\ & ( !\vAluSrc2~0_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_vAluSrc2~0_combout\,
	datae => \ALT_INV_R.aluOp.ALUOpSLTU~q\,
	dataf => \ALT_INV_Mux20~1_combout\,
	combout => \R.aluOp.ALUOpSLTU_OTERM571\);

-- Location: FF_X75_Y5_N44
\R.aluOp.ALUOpSLTU\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \R.aluOp.ALUOpSLTU_OTERM571\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluOp.ALUOpSLTU~q\);

-- Location: LABCELL_X81_Y2_N24
\Mux221~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux221~0_combout\ = ( \R.curInst\(13) & ( !\R.curInst\(12) & ( !\R.curInst\(14) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.curInst\(14),
	datae => \ALT_INV_R.curInst\(13),
	dataf => \ALT_INV_R.curInst\(12),
	combout => \Mux221~0_combout\);

-- Location: LABCELL_X80_Y2_N51
\Mux19~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux19~0_combout\ = ( !\R.curInst\(6) & ( (!\R.curInst\(3) & ((!\R.curInst\(2) & (\Mux221~0_combout\ & (\R.curInst\(4)))) # (\R.curInst\(2) & (((!\R.curInst\(4) & \R.aluOp.ALUOpSLT~q\)))))) # (\R.curInst\(3) & ((((\R.aluOp.ALUOpSLT~q\))))) ) ) # ( 
-- \R.curInst\(6) & ( (\R.aluOp.ALUOpSLT~q\ & ((!\R.curInst\(5)) # (((\R.curInst\(3) & !\R.curInst\(2))) # (\R.curInst\(4))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001000000000000000000001110111010111011111010011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(3),
	datab => \ALT_INV_R.curInst\(2),
	datac => \ALT_INV_R.curInst\(5),
	datad => \ALT_INV_R.curInst\(4),
	datae => \ALT_INV_R.curInst\(6),
	dataf => \ALT_INV_R.aluOp.ALUOpSLT~q\,
	datag => \ALT_INV_Mux221~0_combout\,
	combout => \Mux19~0_combout\);

-- Location: LABCELL_X80_Y2_N21
\R.aluOp.ALUOpSLT_NEW572\ : cyclonev_lcell_comb
-- Equation(s):
-- \R.aluOp.ALUOpSLT_OTERM573\ = ( \R.aluOp.ALUOpSLT~q\ & ( \Mux19~0_combout\ ) ) # ( !\R.aluOp.ALUOpSLT~q\ & ( \Mux19~0_combout\ & ( \vAluSrc2~0_combout\ ) ) ) # ( \R.aluOp.ALUOpSLT~q\ & ( !\Mux19~0_combout\ & ( !\vAluSrc2~0_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101001010101010101011111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_vAluSrc2~0_combout\,
	datae => \ALT_INV_R.aluOp.ALUOpSLT~q\,
	dataf => \ALT_INV_Mux19~0_combout\,
	combout => \R.aluOp.ALUOpSLT_OTERM573\);

-- Location: FF_X80_Y2_N22
\R.aluOp.ALUOpSLT\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \R.aluOp.ALUOpSLT_OTERM573\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluOp.ALUOpSLT~q\);

-- Location: LABCELL_X85_Y5_N24
\Selector32~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector32~0_combout\ = ( !\R.aluOp.ALUOpSLT~q\ & ( !\R.aluOp.ALUOpSLTU~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1100110011001100110011001100110000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluOp.ALUOpSLTU~q\,
	dataf => \ALT_INV_R.aluOp.ALUOpSLT~q\,
	combout => \Selector32~0_combout\);

-- Location: LABCELL_X80_Y5_N0
\LessThan1~32\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~32_combout\ = ( !\LessThan1~28_OTERM51\ & ( !\LessThan1~31_combout\ & ( (!\LessThan1~29_OTERM47\ & (!\LessThan1~30_OTERM43\ & (!\R.aluData1\(25) $ (\R.aluData2\(25))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000010000000000000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData1\(25),
	datab => \ALT_INV_LessThan1~29_OTERM47\,
	datac => \ALT_INV_R.aluData2\(25),
	datad => \ALT_INV_LessThan1~30_OTERM43\,
	datae => \ALT_INV_LessThan1~28_OTERM51\,
	dataf => \ALT_INV_LessThan1~31_combout\,
	combout => \LessThan1~32_combout\);

-- Location: LABCELL_X74_Y5_N57
\LessThan1~0_RTM0345\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~0_RTM0345_combout\ = ( \NxR.aluData2[20]~1_combout\ & ( (!\Mux234~0_combout\) # (!\Mux233~0_combout\ $ (!\NxR.aluData2[21]~0_combout\)) ) ) # ( !\NxR.aluData2[20]~1_combout\ & ( (!\Mux233~0_combout\ $ (!\NxR.aluData2[21]~0_combout\)) # 
-- (\Mux234~0_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101111110101111010111111010111111110101111110101111010111111010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux233~0_combout\,
	datac => \ALT_INV_Mux234~0_combout\,
	datad => \ALT_INV_NxR.aluData2[21]~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[20]~1_combout\,
	combout => \LessThan1~0_RTM0345_combout\);

-- Location: FF_X74_Y5_N58
\LessThan1~0_NEW_REG342\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \LessThan1~0_RTM0345_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \LessThan1~0_OTERM343\);

-- Location: MLABCELL_X72_Y5_N0
\LessThan1~2_RTM0333\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~2_RTM0333_combout\ = ( \Mux237~0_combout\ & ( (!\NxR.aluData2[17]~4_combout\) # (!\NxR.aluData2[16]~5_combout\ $ (!\Mux238~0_combout\)) ) ) # ( !\Mux237~0_combout\ & ( (!\NxR.aluData2[16]~5_combout\ $ (!\Mux238~0_combout\)) # 
-- (\NxR.aluData2[17]~4_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101101011111111010110101111111111111111010110101111111101011010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_NxR.aluData2[16]~5_combout\,
	datac => \ALT_INV_Mux238~0_combout\,
	datad => \ALT_INV_NxR.aluData2[17]~4_combout\,
	dataf => \ALT_INV_Mux237~0_combout\,
	combout => \LessThan1~2_RTM0333_combout\);

-- Location: FF_X72_Y5_N2
\LessThan1~2_NEW_REG330\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \LessThan1~2_RTM0333_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \LessThan1~2_OTERM331\);

-- Location: LABCELL_X75_Y4_N12
\LessThan1~1_RTM0339\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~1_RTM0339_combout\ = ( \NxR.aluData2[18]~3_combout\ & ( (!\Mux236~0_combout\) # (!\NxR.aluData2[19]~2_combout\ $ (!\Mux235~0_combout\)) ) ) # ( !\NxR.aluData2[18]~3_combout\ & ( (!\NxR.aluData2[19]~2_combout\ $ (!\Mux235~0_combout\)) # 
-- (\Mux236~0_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011110011111111001111001111111111111111001111001111111100111100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_NxR.aluData2[19]~2_combout\,
	datac => \ALT_INV_Mux235~0_combout\,
	datad => \ALT_INV_Mux236~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[18]~3_combout\,
	combout => \LessThan1~1_RTM0339_combout\);

-- Location: FF_X75_Y4_N13
\LessThan1~1_NEW_REG336\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \LessThan1~1_RTM0339_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \LessThan1~1_OTERM337\);

-- Location: LABCELL_X75_Y6_N30
\LessThan1~3_RTM0327\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~3_RTM0327_combout\ = ( \NxR.aluData2[15]~6_combout\ & ( (!\Mux239~0_combout\) # (!\NxR.aluData2[14]~7_combout\ $ (!\Mux240~0_combout\)) ) ) # ( !\NxR.aluData2[15]~6_combout\ & ( (!\NxR.aluData2[14]~7_combout\ $ (!\Mux240~0_combout\)) # 
-- (\Mux239~0_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011111111110011001111111111001111001111111111001100111111111100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Mux239~0_combout\,
	datac => \ALT_INV_NxR.aluData2[14]~7_combout\,
	datad => \ALT_INV_Mux240~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[15]~6_combout\,
	combout => \LessThan1~3_RTM0327_combout\);

-- Location: FF_X75_Y6_N32
\LessThan1~3_NEW_REG324\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \LessThan1~3_RTM0327_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \LessThan1~3_OTERM325\);

-- Location: LABCELL_X71_Y6_N12
\LessThan1~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~25_combout\ = ( \Mux241~0_combout\ & ( \NxR.aluData2[13]~10_combout\ & ( (!\Mux242~0_combout\ & \NxR.aluData2[12]~11_combout\) ) ) ) # ( !\Mux241~0_combout\ & ( \NxR.aluData2[13]~10_combout\ ) ) # ( !\Mux241~0_combout\ & ( 
-- !\NxR.aluData2[13]~10_combout\ & ( (!\Mux242~0_combout\ & \NxR.aluData2[12]~11_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011001100000000000000000011111111111111110000000011001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Mux242~0_combout\,
	datad => \ALT_INV_NxR.aluData2[12]~11_combout\,
	datae => \ALT_INV_Mux241~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[13]~10_combout\,
	combout => \LessThan1~25_combout\);

-- Location: FF_X71_Y6_N13
\LessThan1~25_NEW_REG316\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \LessThan1~25_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \LessThan1~25_OTERM317\);

-- Location: LABCELL_X75_Y6_N24
\LessThan1~24\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~24_combout\ = ( \NxR.aluData2[15]~6_combout\ & ( (!\Mux239~0_combout\) # ((!\Mux240~0_combout\ & \NxR.aluData2[14]~7_combout\)) ) ) # ( !\NxR.aluData2[15]~6_combout\ & ( (!\Mux240~0_combout\ & (\NxR.aluData2[14]~7_combout\ & 
-- !\Mux239~0_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101000000000000010100000000011111111000010101111111100001010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux240~0_combout\,
	datac => \ALT_INV_NxR.aluData2[14]~7_combout\,
	datad => \ALT_INV_Mux239~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[15]~6_combout\,
	combout => \LessThan1~24_combout\);

-- Location: FF_X75_Y6_N26
\LessThan1~24_NEW_REG328\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \LessThan1~24_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \LessThan1~24_OTERM329\);

-- Location: LABCELL_X75_Y6_N36
\LessThan1~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~26_combout\ = ( \LessThan1~25_OTERM317\ & ( \LessThan1~24_OTERM329\ & ( (!\LessThan1~0_OTERM343\ & (!\LessThan1~2_OTERM331\ & !\LessThan1~1_OTERM337\)) ) ) ) # ( !\LessThan1~25_OTERM317\ & ( \LessThan1~24_OTERM329\ & ( (!\LessThan1~0_OTERM343\ 
-- & (!\LessThan1~2_OTERM331\ & !\LessThan1~1_OTERM337\)) ) ) ) # ( \LessThan1~25_OTERM317\ & ( !\LessThan1~24_OTERM329\ & ( (!\LessThan1~0_OTERM343\ & (!\LessThan1~2_OTERM331\ & (!\LessThan1~1_OTERM337\ & !\LessThan1~3_OTERM325\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000100000000000000010000000100000001000000010000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_LessThan1~0_OTERM343\,
	datab => \ALT_INV_LessThan1~2_OTERM331\,
	datac => \ALT_INV_LessThan1~1_OTERM337\,
	datad => \ALT_INV_LessThan1~3_OTERM325\,
	datae => \ALT_INV_LessThan1~25_OTERM317\,
	dataf => \ALT_INV_LessThan1~24_OTERM329\,
	combout => \LessThan1~26_combout\);

-- Location: LABCELL_X75_Y6_N3
\LessThan1~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~4_combout\ = ( \Mux243~0_combout\ & ( (\NxR.aluData2[11]~8_combout\ & (!\Mux244~0_combout\ & \NxR.aluData2[10]~9_combout\)) ) ) # ( !\Mux243~0_combout\ & ( ((!\Mux244~0_combout\ & \NxR.aluData2[10]~9_combout\)) # (\NxR.aluData2[11]~8_combout\) 
-- ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001111110011001100111111001100000000001100000000000000110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_NxR.aluData2[11]~8_combout\,
	datac => \ALT_INV_Mux244~0_combout\,
	datad => \ALT_INV_NxR.aluData2[10]~9_combout\,
	dataf => \ALT_INV_Mux243~0_combout\,
	combout => \LessThan1~4_combout\);

-- Location: FF_X75_Y6_N5
\LessThan1~4_NEW_REG318\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \LessThan1~4_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \LessThan1~4_OTERM319\);

-- Location: LABCELL_X71_Y6_N54
\LessThan1~5_RTM0315\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~5_RTM0315_combout\ = ( \NxR.aluData2[12]~11_combout\ & ( (!\Mux242~0_combout\) # (!\NxR.aluData2[13]~10_combout\ $ (!\Mux241~0_combout\)) ) ) # ( !\NxR.aluData2[12]~11_combout\ & ( (!\NxR.aluData2[13]~10_combout\ $ (!\Mux241~0_combout\)) # 
-- (\Mux242~0_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011110011111111001111001111111111111111001111001111111100111100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_NxR.aluData2[13]~10_combout\,
	datac => \ALT_INV_Mux241~0_combout\,
	datad => \ALT_INV_Mux242~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[12]~11_combout\,
	combout => \LessThan1~5_RTM0315_combout\);

-- Location: FF_X71_Y6_N56
\LessThan1~5_NEW_REG312\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \LessThan1~5_RTM0315_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \LessThan1~5_OTERM313\);

-- Location: LABCELL_X75_Y6_N42
\LessThan1~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~6_combout\ = ( !\LessThan1~1_OTERM337\ & ( !\LessThan1~0_OTERM343\ & ( (\LessThan1~4_OTERM319\ & (!\LessThan1~3_OTERM325\ & (!\LessThan1~5_OTERM313\ & !\LessThan1~2_OTERM331\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100000000000000000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_LessThan1~4_OTERM319\,
	datab => \ALT_INV_LessThan1~3_OTERM325\,
	datac => \ALT_INV_LessThan1~5_OTERM313\,
	datad => \ALT_INV_LessThan1~2_OTERM331\,
	datae => \ALT_INV_LessThan1~1_OTERM337\,
	dataf => \ALT_INV_LessThan1~0_OTERM343\,
	combout => \LessThan1~6_combout\);

-- Location: LABCELL_X75_Y4_N30
\LessThan1~20\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~20_combout\ = ( \NxR.aluData2[18]~3_combout\ & ( (!\NxR.aluData2[19]~2_combout\ & (!\Mux235~0_combout\ & !\Mux236~0_combout\)) # (\NxR.aluData2[19]~2_combout\ & ((!\Mux235~0_combout\) # (!\Mux236~0_combout\))) ) ) # ( 
-- !\NxR.aluData2[18]~3_combout\ & ( (\NxR.aluData2[19]~2_combout\ & !\Mux235~0_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011000000110000001100000011000011110011001100001111001100110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_NxR.aluData2[19]~2_combout\,
	datac => \ALT_INV_Mux235~0_combout\,
	datad => \ALT_INV_Mux236~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[18]~3_combout\,
	combout => \LessThan1~20_combout\);

-- Location: FF_X75_Y4_N31
\LessThan1~20_NEW_REG340\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \LessThan1~20_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \LessThan1~20_OTERM341\);

-- Location: LABCELL_X74_Y5_N39
\LessThan1~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~22_combout\ = ( \NxR.aluData2[20]~1_combout\ & ( (!\Mux233~0_combout\ & ((!\Mux234~0_combout\) # (\NxR.aluData2[21]~0_combout\))) # (\Mux233~0_combout\ & (!\Mux234~0_combout\ & \NxR.aluData2[21]~0_combout\)) ) ) # ( 
-- !\NxR.aluData2[20]~1_combout\ & ( (!\Mux233~0_combout\ & \NxR.aluData2[21]~0_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000010101010000000001010101010100000111110101010000011111010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux233~0_combout\,
	datac => \ALT_INV_Mux234~0_combout\,
	datad => \ALT_INV_NxR.aluData2[21]~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[20]~1_combout\,
	combout => \LessThan1~22_combout\);

-- Location: FF_X74_Y5_N40
\LessThan1~22_NEW_REG346\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \LessThan1~22_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \LessThan1~22_OTERM347\);

-- Location: MLABCELL_X72_Y5_N54
\LessThan1~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~21_combout\ = ( \NxR.aluData2[16]~5_combout\ & ( (!\Mux238~0_combout\ & ((!\Mux237~0_combout\) # (\NxR.aluData2[17]~4_combout\))) # (\Mux238~0_combout\ & (!\Mux237~0_combout\ & \NxR.aluData2[17]~4_combout\)) ) ) # ( 
-- !\NxR.aluData2[16]~5_combout\ & ( (!\Mux237~0_combout\ & \NxR.aluData2[17]~4_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011110000000000001111000010100000111110101010000011111010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux238~0_combout\,
	datac => \ALT_INV_Mux237~0_combout\,
	datad => \ALT_INV_NxR.aluData2[17]~4_combout\,
	dataf => \ALT_INV_NxR.aluData2[16]~5_combout\,
	combout => \LessThan1~21_combout\);

-- Location: FF_X72_Y5_N55
\LessThan1~21_NEW_REG334\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \LessThan1~21_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \LessThan1~21_OTERM335\);

-- Location: MLABCELL_X72_Y4_N30
\LessThan1~23\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~23_combout\ = ( !\LessThan1~22_OTERM347\ & ( \LessThan1~21_OTERM335\ & ( ((!\LessThan1~20_OTERM341\ & \LessThan1~1_OTERM337\)) # (\LessThan1~0_OTERM343\) ) ) ) # ( !\LessThan1~22_OTERM347\ & ( !\LessThan1~21_OTERM335\ & ( 
-- (!\LessThan1~20_OTERM341\) # (\LessThan1~0_OTERM343\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1011101110111011000000000000000000111011001110110000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_LessThan1~20_OTERM341\,
	datab => \ALT_INV_LessThan1~0_OTERM343\,
	datac => \ALT_INV_LessThan1~1_OTERM337\,
	datae => \ALT_INV_LessThan1~22_OTERM347\,
	dataf => \ALT_INV_LessThan1~21_OTERM335\,
	combout => \LessThan1~23_combout\);

-- Location: LABCELL_X75_Y6_N15
\LessThan1~18_RTM0323\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~18_RTM0323_combout\ = ( \Mux243~0_combout\ & ( (!\NxR.aluData2[11]~8_combout\) # (!\Mux244~0_combout\ $ (!\NxR.aluData2[10]~9_combout\)) ) ) # ( !\Mux243~0_combout\ & ( (!\Mux244~0_combout\ $ (!\NxR.aluData2[10]~9_combout\)) # 
-- (\NxR.aluData2[11]~8_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011111111110011001111111111001111001111111111001100111111111100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_NxR.aluData2[11]~8_combout\,
	datac => \ALT_INV_Mux244~0_combout\,
	datad => \ALT_INV_NxR.aluData2[10]~9_combout\,
	dataf => \ALT_INV_Mux243~0_combout\,
	combout => \LessThan1~18_RTM0323_combout\);

-- Location: FF_X75_Y6_N17
\LessThan1~18_NEW_REG320\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \LessThan1~18_RTM0323_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \LessThan1~18_OTERM321\);

-- Location: LABCELL_X75_Y6_N6
\LessThan1~19\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~19_combout\ = ( !\LessThan1~5_OTERM313\ & ( !\LessThan1~3_OTERM325\ & ( (!\LessThan1~1_OTERM337\ & (!\LessThan1~18_OTERM321\ & (!\LessThan1~0_OTERM343\ & !\LessThan1~2_OTERM331\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000000000000000000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_LessThan1~1_OTERM337\,
	datab => \ALT_INV_LessThan1~18_OTERM321\,
	datac => \ALT_INV_LessThan1~0_OTERM343\,
	datad => \ALT_INV_LessThan1~2_OTERM331\,
	datae => \ALT_INV_LessThan1~5_OTERM313\,
	dataf => \ALT_INV_LessThan1~3_OTERM325\,
	combout => \LessThan1~19_combout\);

-- Location: LABCELL_X74_Y7_N36
\LessThan1~7_RTM0309\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~7_RTM0309_combout\ = ( \NxR.aluData2[8]~13_combout\ & ( (!\Mux246~0_combout\) # (!\Mux245~0_combout\ $ (!\NxR.aluData2[9]~12_combout\)) ) ) # ( !\NxR.aluData2[8]~13_combout\ & ( (!\Mux245~0_combout\ $ (!\NxR.aluData2[9]~12_combout\)) # 
-- (\Mux246~0_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011111111001111001111111100111111110011111111001111001111111100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Mux245~0_combout\,
	datac => \ALT_INV_Mux246~0_combout\,
	datad => \ALT_INV_NxR.aluData2[9]~12_combout\,
	dataf => \ALT_INV_NxR.aluData2[8]~13_combout\,
	combout => \LessThan1~7_RTM0309_combout\);

-- Location: FF_X74_Y7_N37
\LessThan1~7_NEW_REG306\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \LessThan1~7_RTM0309_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \LessThan1~7_OTERM307\);

-- Location: MLABCELL_X72_Y7_N57
\LessThan1~10_RTM0215\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~10_RTM0215_combout\ = ( \NxR.aluData2[3]~18_combout\ & ( (!\Mux251~0_combout\) # (!\Mux252~0_combout\ $ (!\NxR.aluData2[2]~19_combout\)) ) ) # ( !\NxR.aluData2[3]~18_combout\ & ( (!\Mux252~0_combout\ $ (!\NxR.aluData2[2]~19_combout\)) # 
-- (\Mux251~0_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101111111110101010111111111010110101111111110101010111111111010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux251~0_combout\,
	datac => \ALT_INV_Mux252~0_combout\,
	datad => \ALT_INV_NxR.aluData2[2]~19_combout\,
	dataf => \ALT_INV_NxR.aluData2[3]~18_combout\,
	combout => \LessThan1~10_RTM0215_combout\);

-- Location: FF_X72_Y7_N58
\LessThan1~10_NEW_REG212\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \LessThan1~10_RTM0215_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \LessThan1~10_OTERM213\);

-- Location: LABCELL_X74_Y7_N9
\LessThan1~8_RTM0303\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~8_RTM0303_combout\ = ( \NxR.aluData2[7]~14_combout\ & ( (!\Mux247~0_combout\) # (!\Mux248~0_combout\ $ (!\NxR.aluData2[6]~15_combout\)) ) ) # ( !\NxR.aluData2[7]~14_combout\ & ( (!\Mux248~0_combout\ $ (!\NxR.aluData2[6]~15_combout\)) # 
-- (\Mux247~0_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101101011111111010110101111111111111111010110101111111101011010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux248~0_combout\,
	datac => \ALT_INV_NxR.aluData2[6]~15_combout\,
	datad => \ALT_INV_Mux247~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[7]~14_combout\,
	combout => \LessThan1~8_RTM0303_combout\);

-- Location: FF_X74_Y7_N10
\LessThan1~8_NEW_REG300\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \LessThan1~8_RTM0303_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \LessThan1~8_OTERM301\);

-- Location: MLABCELL_X72_Y7_N12
\LessThan1~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~9_combout\ = ( \NxR.aluData2[1]~17_combout\ & ( (!\Mux253~0_combout\) # ((!\Mux254~0_combout\ & \NxR.aluData2[0]~16_combout\)) ) ) # ( !\NxR.aluData2[1]~17_combout\ & ( (!\Mux253~0_combout\ & (!\Mux254~0_combout\ & 
-- \NxR.aluData2[0]~16_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000010100000000000001010000010101010111110101010101011111010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux253~0_combout\,
	datac => \ALT_INV_Mux254~0_combout\,
	datad => \ALT_INV_NxR.aluData2[0]~16_combout\,
	dataf => \ALT_INV_NxR.aluData2[1]~17_combout\,
	combout => \LessThan1~9_combout\);

-- Location: FF_X72_Y7_N13
\LessThan1~9_NEW_REG252\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \LessThan1~9_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \LessThan1~9_OTERM253\);

-- Location: MLABCELL_X72_Y7_N21
\LessThan1~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~11_combout\ = ( \NxR.aluData2[3]~18_combout\ & ( (!\Mux251~0_combout\) # ((!\Mux252~0_combout\ & \NxR.aluData2[2]~19_combout\)) ) ) # ( !\NxR.aluData2[3]~18_combout\ & ( (!\Mux251~0_combout\ & (!\Mux252~0_combout\ & 
-- \NxR.aluData2[2]~19_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000010100000000000001010000010101010111110101010101011111010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux251~0_combout\,
	datac => \ALT_INV_Mux252~0_combout\,
	datad => \ALT_INV_NxR.aluData2[2]~19_combout\,
	dataf => \ALT_INV_NxR.aluData2[3]~18_combout\,
	combout => \LessThan1~11_combout\);

-- Location: FF_X72_Y7_N22
\LessThan1~11_NEW_REG216\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \LessThan1~11_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \LessThan1~11_OTERM217\);

-- Location: MLABCELL_X72_Y5_N42
\LessThan1~12_RTM0193\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~12_RTM0193_combout\ = ( \NxR.aluData2[5]~21_combout\ & ( (!\Mux249~0_combout\) # (!\NxR.aluData2[4]~20_combout\ $ (!\Mux250~0_combout\)) ) ) # ( !\NxR.aluData2[5]~21_combout\ & ( (!\NxR.aluData2[4]~20_combout\ $ (!\Mux250~0_combout\)) # 
-- (\Mux249~0_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101101011111111010110101111111111111111010110101111111101011010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_NxR.aluData2[4]~20_combout\,
	datac => \ALT_INV_Mux250~0_combout\,
	datad => \ALT_INV_Mux249~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[5]~21_combout\,
	combout => \LessThan1~12_RTM0193_combout\);

-- Location: FF_X72_Y5_N43
\LessThan1~12_NEW_REG190\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \LessThan1~12_RTM0193_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \LessThan1~12_OTERM191\);

-- Location: MLABCELL_X72_Y9_N0
\LessThan1~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~13_combout\ = ( \LessThan1~11_OTERM217\ & ( !\LessThan1~12_OTERM191\ & ( (!\LessThan1~7_OTERM307\ & !\LessThan1~8_OTERM301\) ) ) ) # ( !\LessThan1~11_OTERM217\ & ( !\LessThan1~12_OTERM191\ & ( (!\LessThan1~7_OTERM307\ & 
-- (!\LessThan1~10_OTERM213\ & (!\LessThan1~8_OTERM301\ & \LessThan1~9_OTERM253\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000010000000101000001010000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_LessThan1~7_OTERM307\,
	datab => \ALT_INV_LessThan1~10_OTERM213\,
	datac => \ALT_INV_LessThan1~8_OTERM301\,
	datad => \ALT_INV_LessThan1~9_OTERM253\,
	datae => \ALT_INV_LessThan1~11_OTERM217\,
	dataf => \ALT_INV_LessThan1~12_OTERM191\,
	combout => \LessThan1~13_combout\);

-- Location: LABCELL_X74_Y7_N24
\LessThan1~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~14_combout\ = ( \NxR.aluData2[7]~14_combout\ & ( (!\Mux247~0_combout\) # ((\NxR.aluData2[6]~15_combout\ & !\Mux248~0_combout\)) ) ) # ( !\NxR.aluData2[7]~14_combout\ & ( (\NxR.aluData2[6]~15_combout\ & (!\Mux248~0_combout\ & 
-- !\Mux247~0_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011000000000000001100000000000011111111001100001111111100110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_NxR.aluData2[6]~15_combout\,
	datac => \ALT_INV_Mux248~0_combout\,
	datad => \ALT_INV_Mux247~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[7]~14_combout\,
	combout => \LessThan1~14_combout\);

-- Location: FF_X74_Y7_N25
\LessThan1~14_NEW_REG304\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \LessThan1~14_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \LessThan1~14_OTERM305\);

-- Location: LABCELL_X73_Y5_N57
\LessThan1~15\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~15_combout\ = ( \Mux249~0_combout\ & ( (\NxR.aluData2[4]~20_combout\ & (!\Mux250~0_combout\ & \NxR.aluData2[5]~21_combout\)) ) ) # ( !\Mux249~0_combout\ & ( ((\NxR.aluData2[4]~20_combout\ & !\Mux250~0_combout\)) # (\NxR.aluData2[5]~21_combout\) 
-- ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101000011111111010100001111111100000000010100000000000001010000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_NxR.aluData2[4]~20_combout\,
	datac => \ALT_INV_Mux250~0_combout\,
	datad => \ALT_INV_NxR.aluData2[5]~21_combout\,
	dataf => \ALT_INV_Mux249~0_combout\,
	combout => \LessThan1~15_combout\);

-- Location: FF_X73_Y5_N58
\LessThan1~15_NEW_REG194\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \LessThan1~15_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \LessThan1~15_OTERM195\);

-- Location: LABCELL_X74_Y7_N42
\LessThan1~16\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~16_combout\ = ( \NxR.aluData2[8]~13_combout\ & ( (!\Mux245~0_combout\ & ((!\Mux246~0_combout\) # (\NxR.aluData2[9]~12_combout\))) # (\Mux245~0_combout\ & (!\Mux246~0_combout\ & \NxR.aluData2[9]~12_combout\)) ) ) # ( 
-- !\NxR.aluData2[8]~13_combout\ & ( (!\Mux245~0_combout\ & \NxR.aluData2[9]~12_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011001100000000001100110011000000111111001100000011111100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Mux245~0_combout\,
	datac => \ALT_INV_Mux246~0_combout\,
	datad => \ALT_INV_NxR.aluData2[9]~12_combout\,
	dataf => \ALT_INV_NxR.aluData2[8]~13_combout\,
	combout => \LessThan1~16_combout\);

-- Location: FF_X74_Y7_N44
\LessThan1~16_NEW_REG310\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \LessThan1~16_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \LessThan1~16_OTERM311\);

-- Location: MLABCELL_X72_Y9_N6
\LessThan1~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~17_combout\ = ( \LessThan1~7_OTERM307\ & ( !\LessThan1~16_OTERM311\ ) ) # ( !\LessThan1~7_OTERM307\ & ( !\LessThan1~16_OTERM311\ & ( (!\LessThan1~14_OTERM305\ & ((!\LessThan1~15_OTERM195\) # (\LessThan1~8_OTERM301\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1100010011000100111111111111111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_LessThan1~8_OTERM301\,
	datab => \ALT_INV_LessThan1~14_OTERM305\,
	datac => \ALT_INV_LessThan1~15_OTERM195\,
	datae => \ALT_INV_LessThan1~7_OTERM307\,
	dataf => \ALT_INV_LessThan1~16_OTERM311\,
	combout => \LessThan1~17_combout\);

-- Location: LABCELL_X75_Y6_N18
\LessThan1~27\ : cyclonev_lcell_comb
-- Equation(s):
-- \LessThan1~27_combout\ = ( \LessThan1~13_combout\ & ( \LessThan1~17_combout\ & ( (!\LessThan1~26_combout\ & (!\LessThan1~6_combout\ & (\LessThan1~23_combout\ & !\LessThan1~19_combout\))) ) ) ) # ( !\LessThan1~13_combout\ & ( \LessThan1~17_combout\ & ( 
-- (!\LessThan1~26_combout\ & (!\LessThan1~6_combout\ & \LessThan1~23_combout\)) ) ) ) # ( \LessThan1~13_combout\ & ( !\LessThan1~17_combout\ & ( (!\LessThan1~26_combout\ & (!\LessThan1~6_combout\ & (\LessThan1~23_combout\ & !\LessThan1~19_combout\))) ) ) ) 
-- # ( !\LessThan1~13_combout\ & ( !\LessThan1~17_combout\ & ( (!\LessThan1~26_combout\ & (!\LessThan1~6_combout\ & (\LessThan1~23_combout\ & !\LessThan1~19_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000100000000000000010000000000000001000000010000000100000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_LessThan1~26_combout\,
	datab => \ALT_INV_LessThan1~6_combout\,
	datac => \ALT_INV_LessThan1~23_combout\,
	datad => \ALT_INV_LessThan1~19_combout\,
	datae => \ALT_INV_LessThan1~13_combout\,
	dataf => \ALT_INV_LessThan1~17_combout\,
	combout => \LessThan1~27_combout\);

-- Location: LABCELL_X80_Y5_N42
\Selector32~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector32~1_combout\ = ( \LessThan1~32_combout\ & ( \LessThan1~27_combout\ & ( (!\Selector32~0_combout\ & (((!\LessThan1~36_combout\ & \LessThan1~37_combout\)) # (\LessThan1~38_combout\))) ) ) ) # ( !\LessThan1~32_combout\ & ( \LessThan1~27_combout\ & ( 
-- (!\Selector32~0_combout\ & (((!\LessThan1~36_combout\ & \LessThan1~37_combout\)) # (\LessThan1~38_combout\))) ) ) ) # ( \LessThan1~32_combout\ & ( !\LessThan1~27_combout\ & ( (!\Selector32~0_combout\ & ((\LessThan1~37_combout\) # 
-- (\LessThan1~38_combout\))) ) ) ) # ( !\LessThan1~32_combout\ & ( !\LessThan1~27_combout\ & ( (!\Selector32~0_combout\ & (((!\LessThan1~36_combout\ & \LessThan1~37_combout\)) # (\LessThan1~38_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011101100000000001111110000000000111011000000000011101100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_LessThan1~36_combout\,
	datab => \ALT_INV_LessThan1~38_combout\,
	datac => \ALT_INV_LessThan1~37_combout\,
	datad => \ALT_INV_Selector32~0_combout\,
	datae => \ALT_INV_LessThan1~32_combout\,
	dataf => \ALT_INV_LessThan1~27_combout\,
	combout => \Selector32~1_combout\);

-- Location: LABCELL_X80_Y5_N21
\Selector32~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector32~8_combout\ = ( \Selector32~1_combout\ ) # ( !\Selector32~1_combout\ & ( !\Selector32~7_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010101010101010101010101010101011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector32~7_combout\,
	dataf => \ALT_INV_Selector32~1_combout\,
	combout => \Selector32~8_combout\);

-- Location: FF_X80_Y5_N23
\R.aluRes[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector32~8_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.aluCalc~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluRes\(0));

-- Location: LABCELL_X80_Y5_N12
\Comb:vRegWriteData[0]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vRegWriteData[0]~1_combout\ = ( \R.aluRes\(0) & ( \Selector32~1_combout\ & ( (!\R.memToReg~q\) # (\Comb:vRegWriteData[0]~0_combout\) ) ) ) # ( !\R.aluRes\(0) & ( \Selector32~1_combout\ & ( ((\R.aluCalc~q\ & !\R.memToReg~q\)) # 
-- (\Comb:vRegWriteData[0]~0_combout\) ) ) ) # ( \R.aluRes\(0) & ( !\Selector32~1_combout\ & ( ((!\R.memToReg~q\ & ((!\Selector32~7_combout\) # (!\R.aluCalc~q\)))) # (\Comb:vRegWriteData[0]~0_combout\) ) ) ) # ( !\R.aluRes\(0) & ( !\Selector32~1_combout\ & ( 
-- ((!\Selector32~7_combout\ & (\R.aluCalc~q\ & !\R.memToReg~q\))) # (\Comb:vRegWriteData[0]~0_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011101100110011111110110011001100111111001100111111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector32~7_combout\,
	datab => \ALT_INV_Comb:vRegWriteData[0]~0_combout\,
	datac => \ALT_INV_R.aluCalc~q\,
	datad => \ALT_INV_R.memToReg~q\,
	datae => \ALT_INV_R.aluRes\(0),
	dataf => \ALT_INV_Selector32~1_combout\,
	combout => \Comb:vRegWriteData[0]~1_combout\);

-- Location: FF_X80_Y5_N8
\R.curPC[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[0]~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC\(0));

-- Location: FF_X80_Y5_N14
\R.regWriteData[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vRegWriteData[0]~1_combout\,
	asdata => \R.curPC\(0),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.regWriteData\(0));

-- Location: FF_X72_Y6_N26
\RegFile[3][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(0),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~6_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[3][0]~q\);

-- Location: LABCELL_X68_Y6_N6
\Mux122~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux122~0_combout\ = ( \R.curInst\(21) & ( \R.curInst\(20) & ( \RegFile[7][0]~q\ ) ) ) # ( !\R.curInst\(21) & ( \R.curInst\(20) & ( \RegFile[5][0]~q\ ) ) ) # ( \R.curInst\(21) & ( !\R.curInst\(20) & ( \RegFile[6][0]~q\ ) ) ) # ( !\R.curInst\(21) & ( 
-- !\R.curInst\(20) & ( \RegFile[4][0]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111001100110011001101010101010101010000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[5][0]~q\,
	datab => \ALT_INV_RegFile[6][0]~q\,
	datac => \ALT_INV_RegFile[7][0]~q\,
	datad => \ALT_INV_RegFile[4][0]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	combout => \Mux122~0_combout\);

-- Location: MLABCELL_X72_Y6_N24
\Mux122~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux122~26_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((\RegFile[1][0]~q\ & (\R.curInst\(20)))))) # (\R.curInst\(22) & ((((\Mux122~0_combout\))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & ((!\R.curInst\(20) & (((\RegFile[2][0]~q\)))) # 
-- (\R.curInst\(20) & (\RegFile[3][0]~q\)))) # (\R.curInst\(22) & ((((\Mux122~0_combout\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001010000010100010001001010101010111110101111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(22),
	datab => \ALT_INV_RegFile[3][0]~q\,
	datac => \ALT_INV_RegFile[2][0]~q\,
	datad => \ALT_INV_R.curInst\(20),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux122~0_combout\,
	datag => \ALT_INV_RegFile[1][0]~q\,
	combout => \Mux122~26_combout\);

-- Location: MLABCELL_X72_Y6_N30
\Mux122~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux122~22_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & (\RegFile[24][0]~q\)) # (\R.curInst\(20) & ((\RegFile[25][0]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( (!\R.curInst\(22) & 
-- (((!\R.curInst\(20) & ((\RegFile[26][0]~q\))) # (\R.curInst\(20) & (\RegFile[27][0]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110000110011111111110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[27][0]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[26][0]~q\,
	datad => \ALT_INV_RegFile[25][0]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[24][0]~q\,
	combout => \Mux122~22_combout\);

-- Location: FF_X71_Y8_N32
\RegFile[28][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[28][0]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~17_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[28][0]~q\);

-- Location: MLABCELL_X72_Y6_N42
\Mux122~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux122~9_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux122~22_combout\))))) # (\R.curInst\(22) & (((!\Mux122~22_combout\ & ((\RegFile[28][0]~q\))) # (\Mux122~22_combout\ & (\RegFile[29][0]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux122~22_combout\)))) # (\R.curInst\(22) & ((!\Mux122~22_combout\ & (\RegFile[30][0]~q\)) # (\Mux122~22_combout\ & ((\RegFile[31][0]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[29][0]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[30][0]~q\,
	datad => \ALT_INV_RegFile[31][0]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux122~22_combout\,
	datag => \ALT_INV_RegFile[28][0]~q\,
	combout => \Mux122~9_combout\);

-- Location: FF_X66_Y4_N17
\RegFile[18][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \RegFile[18][0]~feeder_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \Decoder0~26_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[18][0]~q\);

-- Location: LABCELL_X66_Y4_N48
\Mux122~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux122~18_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & ((!\R.curInst\(20) & ((\RegFile[16][0]~q\))) # (\R.curInst\(20) & (\RegFile[17][0]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & ((\RegFile[18][0]~q\))) # (\R.curInst\(20) & (\RegFile[19][0]~q\)))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000111100000000000011110000000000110011111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[19][0]~q\,
	datab => \ALT_INV_RegFile[17][0]~q\,
	datac => \ALT_INV_RegFile[18][0]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[16][0]~q\,
	combout => \Mux122~18_combout\);

-- Location: MLABCELL_X72_Y6_N0
\Mux122~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux122~5_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & ((((\Mux122~18_combout\))))) # (\R.curInst\(22) & (((!\Mux122~18_combout\ & ((\RegFile[20][0]~q\))) # (\Mux122~18_combout\ & (\RegFile[21][0]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux122~18_combout\)))) # (\R.curInst\(22) & ((!\Mux122~18_combout\ & (\RegFile[22][0]~q\)) # (\Mux122~18_combout\ & ((\RegFile[23][0]~q\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000001100000011000000110000001111011101110111011100110011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[21][0]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[22][0]~q\,
	datad => \ALT_INV_RegFile[23][0]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux122~18_combout\,
	datag => \ALT_INV_RegFile[20][0]~q\,
	combout => \Mux122~5_combout\);

-- Location: LABCELL_X66_Y8_N12
\Mux122~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux122~14_combout\ = ( !\R.curInst\(21) & ( (!\R.curInst\(22) & (((!\R.curInst\(20) & ((\RegFile[8][0]~q\))) # (\R.curInst\(20) & (\RegFile[9][0]~q\))))) # (\R.curInst\(22) & ((((\R.curInst\(20)))))) ) ) # ( \R.curInst\(21) & ( ((!\R.curInst\(22) & 
-- ((!\R.curInst\(20) & (\RegFile[10][0]~q\)) # (\R.curInst\(20) & ((\RegFile[11][0]~q\))))) # (\R.curInst\(22) & (((\R.curInst\(20)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000110000001100000011000000110001110111011101110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[9][0]~q\,
	datab => \ALT_INV_R.curInst\(22),
	datac => \ALT_INV_RegFile[10][0]~q\,
	datad => \ALT_INV_RegFile[11][0]~q\,
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_R.curInst\(20),
	datag => \ALT_INV_RegFile[8][0]~q\,
	combout => \Mux122~14_combout\);

-- Location: FF_X70_Y8_N22
\RegFile[12][0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \R.regWriteData\(0),
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \Decoder0~9_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \RegFile[12][0]~q\);

-- Location: LABCELL_X66_Y8_N0
\Mux122~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux122~1_combout\ = ( !\R.curInst\(21) & ( ((!\R.curInst\(22) & (((\Mux122~14_combout\)))) # (\R.curInst\(22) & ((!\Mux122~14_combout\ & ((\RegFile[12][0]~q\))) # (\Mux122~14_combout\ & (\RegFile[13][0]~q\))))) ) ) # ( \R.curInst\(21) & ( 
-- ((!\R.curInst\(22) & (((\Mux122~14_combout\)))) # (\R.curInst\(22) & ((!\Mux122~14_combout\ & ((\RegFile[14][0]~q\))) # (\Mux122~14_combout\ & (\RegFile[15][0]~q\))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000001111000000000000111111111111001100111111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_RegFile[15][0]~q\,
	datab => \ALT_INV_RegFile[13][0]~q\,
	datac => \ALT_INV_RegFile[14][0]~q\,
	datad => \ALT_INV_R.curInst\(22),
	datae => \ALT_INV_R.curInst\(21),
	dataf => \ALT_INV_Mux122~14_combout\,
	datag => \ALT_INV_RegFile[12][0]~q\,
	combout => \Mux122~1_combout\);

-- Location: MLABCELL_X72_Y6_N36
\Mux122~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux122~13_combout\ = ( \Mux122~5_combout\ & ( \Mux122~1_combout\ & ( (!\R.curInst\(24) & (((\Mux122~26_combout\)) # (\R.curInst\(23)))) # (\R.curInst\(24) & ((!\R.curInst\(23)) # ((\Mux122~9_combout\)))) ) ) ) # ( !\Mux122~5_combout\ & ( 
-- \Mux122~1_combout\ & ( (!\R.curInst\(24) & (((\Mux122~26_combout\)) # (\R.curInst\(23)))) # (\R.curInst\(24) & (\R.curInst\(23) & ((\Mux122~9_combout\)))) ) ) ) # ( \Mux122~5_combout\ & ( !\Mux122~1_combout\ & ( (!\R.curInst\(24) & (!\R.curInst\(23) & 
-- (\Mux122~26_combout\))) # (\R.curInst\(24) & ((!\R.curInst\(23)) # ((\Mux122~9_combout\)))) ) ) ) # ( !\Mux122~5_combout\ & ( !\Mux122~1_combout\ & ( (!\R.curInst\(24) & (!\R.curInst\(23) & (\Mux122~26_combout\))) # (\R.curInst\(24) & (\R.curInst\(23) & 
-- ((\Mux122~9_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000100000011001010011000101110100101010001110110110111001111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(24),
	datab => \ALT_INV_R.curInst\(23),
	datac => \ALT_INV_Mux122~26_combout\,
	datad => \ALT_INV_Mux122~9_combout\,
	datae => \ALT_INV_Mux122~5_combout\,
	dataf => \ALT_INV_Mux122~1_combout\,
	combout => \Mux122~13_combout\);

-- Location: LABCELL_X73_Y6_N18
\NxR.aluData2[0]~16\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR.aluData2[0]~16_combout\ = ( \Mux122~13_combout\ & ( (!\vAluSrc2~1_combout\) # ((\Mux154~1_combout\ & (!\R.curInst\(3) & \Equal4~1_combout\))) ) ) # ( !\Mux122~13_combout\ & ( (\Mux154~1_combout\ & (!\R.curInst\(3) & (\vAluSrc2~1_combout\ & 
-- \Equal4~1_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000100000000000000010011110000111101001111000011110100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux154~1_combout\,
	datab => \ALT_INV_R.curInst\(3),
	datac => \ALT_INV_vAluSrc2~1_combout\,
	datad => \ALT_INV_Equal4~1_combout\,
	dataf => \ALT_INV_Mux122~13_combout\,
	combout => \NxR.aluData2[0]~16_combout\);

-- Location: FF_X73_Y6_N46
\R.aluData2[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	asdata => \NxR.aluData2[0]~16_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.aluData2\(0));

-- Location: LABCELL_X71_Y7_N24
\Selector32~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector32~4_combout\ = ( \NxR.aluData2[0]~16_combout\ & ( ((\R.aluOp.ALUOpAnd_OTERM357\ & \Mux254~0_combout\)) # (\R.aluOp.ALUOpOr_OTERM353\) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( (\R.aluOp.ALUOpOr_OTERM353\ & \Mux254~0_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110011000000000011001100110011001111110011001100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluOp.ALUOpOr_OTERM353\,
	datac => \ALT_INV_R.aluOp.ALUOpAnd_OTERM357\,
	datad => \ALT_INV_Mux254~0_combout\,
	dataf => \ALT_INV_NxR.aluData2[0]~16_combout\,
	combout => \Selector32~4_combout\);

-- Location: FF_X71_Y7_N25
\Selector32~4_NEW_REG396\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Selector32~4_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Selector32~4_OTERM397\);

-- Location: LABCELL_X80_Y7_N3
\Selector32~7_RESYN1056\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector32~7_RESYN1056_BDD1057\ = ( \ShiftLeft0~0_OTERM263\ & ( (!\Selector32~3_OTERM379\ & !\Selector32~4_OTERM397\) ) ) # ( !\ShiftLeft0~0_OTERM263\ & ( !\Selector32~4_OTERM397\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111000011110000111100001111000011000000110000001100000011000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Selector32~3_OTERM379\,
	datac => \ALT_INV_Selector32~4_OTERM397\,
	dataf => \ALT_INV_ShiftLeft0~0_OTERM263\,
	combout => \Selector32~7_RESYN1056_BDD1057\);

-- Location: LABCELL_X81_Y7_N36
\Selector32~7_RESYN1058\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector32~7_RESYN1058_BDD1059\ = ( \R.aluData1\(31) & ( (\Selector32~7_RESYN1056_BDD1057\ & ((!\R.aluOp.ALUOpSLT~q\) # (\R.aluData2\(31)))) ) ) # ( !\R.aluData1\(31) & ( (\Selector32~7_RESYN1056_BDD1057\ & ((!\R.aluData2\(31)) # 
-- (!\R.aluOp.ALUOpSLTU~q\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100100010001100110010001000110001001100010011000100110001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(31),
	datab => \ALT_INV_Selector32~7_RESYN1056_BDD1057\,
	datac => \ALT_INV_R.aluOp.ALUOpSLT~q\,
	datad => \ALT_INV_R.aluOp.ALUOpSLTU~q\,
	dataf => \ALT_INV_R.aluData1\(31),
	combout => \Selector32~7_RESYN1058_BDD1059\);

-- Location: MLABCELL_X72_Y7_N36
\ShiftRight1~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~5_combout\ = ( \NxR.aluData2[0]~16_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( \Mux251~0_combout\ ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( \NxR.aluData2[1]~17_combout\ & ( \Mux252~0_combout\ ) ) ) # ( \NxR.aluData2[0]~16_combout\ & ( 
-- !\NxR.aluData2[1]~17_combout\ & ( \Mux253~0_combout\ ) ) ) # ( !\NxR.aluData2[0]~16_combout\ & ( !\NxR.aluData2[1]~17_combout\ & ( \Mux254~0_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101000011110000111100000000111111110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux254~0_combout\,
	datab => \ALT_INV_Mux251~0_combout\,
	datac => \ALT_INV_Mux253~0_combout\,
	datad => \ALT_INV_Mux252~0_combout\,
	datae => \ALT_INV_NxR.aluData2[0]~16_combout\,
	dataf => \ALT_INV_NxR.aluData2[1]~17_combout\,
	combout => \ShiftRight1~5_combout\);

-- Location: FF_X72_Y7_N37
\ShiftRight1~5_NEW_REG218\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \ShiftRight1~5_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ShiftRight1~5_OTERM219\);

-- Location: LABCELL_X74_Y8_N24
\ShiftRight1~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \ShiftRight1~9_combout\ = ( \R.aluData2\(3) & ( \R.aluData2\(2) & ( \ShiftRight1~8_OTERM261\ ) ) ) # ( !\R.aluData2\(3) & ( \R.aluData2\(2) & ( \ShiftRight1~6_OTERM197\ ) ) ) # ( \R.aluData2\(3) & ( !\R.aluData2\(2) & ( \ShiftRight1~7_OTERM259\ ) ) ) # ( 
-- !\R.aluData2\(3) & ( !\R.aluData2\(2) & ( \ShiftRight1~5_OTERM219\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101000000001111111100001111000011110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_ShiftRight1~5_OTERM219\,
	datab => \ALT_INV_ShiftRight1~8_OTERM261\,
	datac => \ALT_INV_ShiftRight1~6_OTERM197\,
	datad => \ALT_INV_ShiftRight1~7_OTERM259\,
	datae => \ALT_INV_R.aluData2\(3),
	dataf => \ALT_INV_R.aluData2\(2),
	combout => \ShiftRight1~9_combout\);

-- Location: LABCELL_X80_Y5_N57
\Selector32~7_RESYN1060\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector32~7_RESYN1060_BDD1061\ = ( \ShiftRight1~4_combout\ & ( (!\R.aluData2\(4) & !\ShiftRight1~9_combout\) ) ) # ( !\ShiftRight1~4_combout\ & ( (!\ShiftRight1~9_combout\) # (\R.aluData2\(4)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111010111110101111101011111010110100000101000001010000010100000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluData2\(4),
	datac => \ALT_INV_ShiftRight1~9_combout\,
	dataf => \ALT_INV_ShiftRight1~4_combout\,
	combout => \Selector32~7_RESYN1060_BDD1061\);

-- Location: LABCELL_X81_Y7_N0
\Selector32~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector32~2_combout\ = ( \R.aluData2\(0) & ( \R.aluOp.ALUOpXor~DUPLICATE_q\ & ( !\Add2~1_OTERM735_OTERM837\ ) ) ) # ( !\R.aluData2\(0) & ( \R.aluOp.ALUOpXor~DUPLICATE_q\ & ( \Add2~1_OTERM735_OTERM837\ ) ) ) # ( \R.aluData2\(0) & ( 
-- !\R.aluOp.ALUOpXor~DUPLICATE_q\ & ( (\R.aluOp.ALUOpAdd~q\ & !\Add2~1_OTERM735_OTERM837\) ) ) ) # ( !\R.aluData2\(0) & ( !\R.aluOp.ALUOpXor~DUPLICATE_q\ & ( (\R.aluOp.ALUOpAdd~q\ & \Add2~1_OTERM735_OTERM837\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011001100000011000000001111000011111111000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datac => \ALT_INV_Add2~1_OTERM735_OTERM837\,
	datae => \ALT_INV_R.aluData2\(0),
	dataf => \ALT_INV_R.aluOp.ALUOpXor~DUPLICATE_q\,
	combout => \Selector32~2_combout\);

-- Location: LABCELL_X80_Y5_N24
\Selector32~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector32~7_combout\ = ( \Selector32~7_RESYN1060_BDD1061\ & ( !\Selector32~2_combout\ & ( (\Selector32~7_RESYN1058_BDD1059\ & ((!\Add2~1_sumout\) # (!\R.aluOp.ALUOpSub~q\))) ) ) ) # ( !\Selector32~7_RESYN1060_BDD1061\ & ( !\Selector32~2_combout\ & ( 
-- (!\Selector31~0_OTERM349\ & (\Selector32~7_RESYN1058_BDD1059\ & ((!\Add2~1_sumout\) # (!\R.aluOp.ALUOpSub~q\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000110000001000000011110000101000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add2~1_sumout\,
	datab => \ALT_INV_Selector31~0_OTERM349\,
	datac => \ALT_INV_Selector32~7_RESYN1058_BDD1059\,
	datad => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datae => \ALT_INV_Selector32~7_RESYN1060_BDD1061\,
	dataf => \ALT_INV_Selector32~2_combout\,
	combout => \Selector32~7_combout\);

-- Location: LABCELL_X80_Y5_N6
\Comb:vJumpAdr[0]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Comb:vJumpAdr[0]~0_combout\ = ( \Add3~1_sumout\ & ( \Selector32~1_combout\ & ( ((!\Equal4~2_combout\) # (\R.aluCalc~q\)) # (\R.aluRes[0]~DUPLICATE_q\) ) ) ) # ( !\Add3~1_sumout\ & ( \Selector32~1_combout\ & ( (\Equal4~2_combout\ & ((\R.aluCalc~q\) # 
-- (\R.aluRes[0]~DUPLICATE_q\))) ) ) ) # ( \Add3~1_sumout\ & ( !\Selector32~1_combout\ & ( (!\Equal4~2_combout\) # ((!\R.aluCalc~q\ & ((\R.aluRes[0]~DUPLICATE_q\))) # (\R.aluCalc~q\ & (!\Selector32~7_combout\))) ) ) ) # ( !\Add3~1_sumout\ & ( 
-- !\Selector32~1_combout\ & ( (\Equal4~2_combout\ & ((!\R.aluCalc~q\ & ((\R.aluRes[0]~DUPLICATE_q\))) # (\R.aluCalc~q\ & (!\Selector32~7_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000111010111111110011101000000000001111111111111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector32~7_combout\,
	datab => \ALT_INV_R.aluRes[0]~DUPLICATE_q\,
	datac => \ALT_INV_R.aluCalc~q\,
	datad => \ALT_INV_Equal4~2_combout\,
	datae => \ALT_INV_Add3~1_sumout\,
	dataf => \ALT_INV_Selector32~1_combout\,
	combout => \Comb:vJumpAdr[0]~0_combout\);

-- Location: FF_X80_Y5_N7
\R.curPC[0]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[0]~0_combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	ena => \R.jumpToAdr~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC[0]~DUPLICATE_q\);

-- Location: FF_X78_Y4_N14
\R.curPC[29]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \Comb:vJumpAdr[29]~0_combout\,
	asdata => \Add0~109_sumout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sload => \ALT_INV_R.jumpToAdr~q\,
	ena => \NxR.curPC[31]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.curPC[29]~DUPLICATE_q\);

-- Location: LABCELL_X80_Y3_N48
\vAluRes~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~9_combout\ = (!\R.aluCalc~q\ & (\R.aluRes\(9))) # (\R.aluCalc~q\ & (((!\Selector23~5_combout\) # (\Selector23~0_combout\))))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0111011100100111011101110010011101110111001001110111011100100111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluCalc~q\,
	datab => \ALT_INV_R.aluRes\(9),
	datac => \ALT_INV_Selector23~0_combout\,
	datad => \ALT_INV_Selector23~5_combout\,
	combout => \vAluRes~9_combout\);

-- Location: LABCELL_X81_Y4_N42
\vAluRes~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~11_combout\ = ( \Selector20~4_combout\ & ( (\R.aluRes\(12)) # (\R.aluCalc~q\) ) ) # ( !\Selector20~4_combout\ & ( (!\R.aluCalc~q\ & ((\R.aluRes\(12)))) # (\R.aluCalc~q\ & (!\Selector20~3_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101011111010000010101111101000001111111111110000111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector20~3_combout\,
	datac => \ALT_INV_R.aluCalc~q\,
	datad => \ALT_INV_R.aluRes\(12),
	dataf => \ALT_INV_Selector20~4_combout\,
	combout => \vAluRes~11_combout\);

-- Location: MLABCELL_X78_Y3_N42
\vAluRes~12\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~12_combout\ = ( \Selector18~3_combout\ & ( (!\R.aluCalc~q\ & (\R.aluRes\(14))) # (\R.aluCalc~q\ & ((\Selector18~4_combout\))) ) ) # ( !\Selector18~3_combout\ & ( (\R.aluRes\(14)) # (\R.aluCalc~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011111100111111001111110011111100001100001111110000110000111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_R.aluRes\(14),
	datad => \ALT_INV_Selector18~4_combout\,
	dataf => \ALT_INV_Selector18~3_combout\,
	combout => \vAluRes~12_combout\);

-- Location: LABCELL_X79_Y3_N27
\Selector16~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector16~4_combout\ = ( \Add2~65_sumout\ & ( ((\R.aluOp.ALUOpAdd~q\ & \Add1~65_sumout\)) # (\R.aluOp.ALUOpSub~q\) ) ) # ( !\Add2~65_sumout\ & ( (\R.aluOp.ALUOpAdd~q\ & \Add1~65_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010101000000000101010100001111010111110000111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	datac => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datad => \ALT_INV_Add1~65_sumout\,
	dataf => \ALT_INV_Add2~65_sumout\,
	combout => \Selector16~4_combout\);

-- Location: LABCELL_X79_Y3_N24
\vAluRes~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~13_combout\ = ( \R.aluRes\(16) & ( (!\R.aluCalc~q\) # ((!\Selector16~3_combout\) # (\Selector16~4_combout\)) ) ) # ( !\R.aluRes\(16) & ( (\R.aluCalc~q\ & ((!\Selector16~3_combout\) # (\Selector16~4_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100000011001100110000001111111111110011111111111111001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_Selector16~4_combout\,
	datad => \ALT_INV_Selector16~3_combout\,
	dataf => \ALT_INV_R.aluRes\(16),
	combout => \vAluRes~13_combout\);

-- Location: MLABCELL_X78_Y3_N48
\Selector15~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Selector15~1_combout\ = ( \Add1~69_sumout\ & ( \R.aluOp.ALUOpAdd~q\ ) ) # ( !\Add1~69_sumout\ & ( \R.aluOp.ALUOpAdd~q\ & ( (\Add2~69_sumout\ & \R.aluOp.ALUOpSub~q\) ) ) ) # ( \Add1~69_sumout\ & ( !\R.aluOp.ALUOpAdd~q\ & ( (\Add2~69_sumout\ & 
-- \R.aluOp.ALUOpSub~q\) ) ) ) # ( !\Add1~69_sumout\ & ( !\R.aluOp.ALUOpAdd~q\ & ( (\Add2~69_sumout\ & \R.aluOp.ALUOpSub~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100010001000100010001000100010001000100011111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Add2~69_sumout\,
	datab => \ALT_INV_R.aluOp.ALUOpSub~q\,
	datae => \ALT_INV_Add1~69_sumout\,
	dataf => \ALT_INV_R.aluOp.ALUOpAdd~q\,
	combout => \Selector15~1_combout\);

-- Location: MLABCELL_X78_Y3_N24
\vAluRes~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~14_combout\ = ( \R.aluRes\(17) & ( \Selector15~4_combout\ & ( ((!\R.aluCalc~q\) # (\Selector15~0_combout\)) # (\Selector15~1_combout\) ) ) ) # ( !\R.aluRes\(17) & ( \Selector15~4_combout\ & ( (\R.aluCalc~q\ & ((\Selector15~0_combout\) # 
-- (\Selector15~1_combout\))) ) ) ) # ( \R.aluRes\(17) & ( !\Selector15~4_combout\ ) ) # ( !\R.aluRes\(17) & ( !\Selector15~4_combout\ & ( \R.aluCalc~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111111111111111111100000000011101111111111101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector15~1_combout\,
	datab => \ALT_INV_Selector15~0_combout\,
	datad => \ALT_INV_R.aluCalc~q\,
	datae => \ALT_INV_R.aluRes\(17),
	dataf => \ALT_INV_Selector15~4_combout\,
	combout => \vAluRes~14_combout\);

-- Location: LABCELL_X79_Y3_N3
\vAluRes~15\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~15_combout\ = ( \R.aluData2\(4) & ( (!\R.aluCalc~q\ & ((\R.aluRes\(18)))) # (\R.aluCalc~q\ & (!\Selector14~3_combout\)) ) ) # ( !\R.aluData2\(4) & ( (!\R.aluCalc~q\ & (((\R.aluRes\(18))))) # (\R.aluCalc~q\ & ((!\Selector14~0_combout\) # 
-- ((!\Selector14~3_combout\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010011111110010101001111111001010000111110100101000011111010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.aluCalc~q\,
	datab => \ALT_INV_Selector14~0_combout\,
	datac => \ALT_INV_Selector14~3_combout\,
	datad => \ALT_INV_R.aluRes\(18),
	dataf => \ALT_INV_R.aluData2\(4),
	combout => \vAluRes~15_combout\);

-- Location: LABCELL_X83_Y4_N57
\vAluRes~16\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~16_combout\ = ( \R.aluCalc~q\ & ( \Selector13~0_combout\ & ( !\Selector13~1_combout\ ) ) ) # ( !\R.aluCalc~q\ & ( \Selector13~0_combout\ & ( \R.aluRes\(19) ) ) ) # ( \R.aluCalc~q\ & ( !\Selector13~0_combout\ & ( (!\Selector13~1_combout\) # 
-- (!\R.aluData2\(4)) ) ) ) # ( !\R.aluCalc~q\ & ( !\Selector13~0_combout\ & ( \R.aluRes\(19) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110011111110101111101000110011001100111010101010101010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Selector13~1_combout\,
	datab => \ALT_INV_R.aluRes\(19),
	datac => \ALT_INV_R.aluData2\(4),
	datae => \ALT_INV_R.aluCalc~q\,
	dataf => \ALT_INV_Selector13~0_combout\,
	combout => \vAluRes~16_combout\);

-- Location: MLABCELL_X78_Y2_N3
\vAluRes~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~18_combout\ = ( \R.aluRes\(21) & ( \R.aluCalc~q\ & ( \Selector11~5_combout\ ) ) ) # ( !\R.aluRes\(21) & ( \R.aluCalc~q\ & ( \Selector11~5_combout\ ) ) ) # ( \R.aluRes\(21) & ( !\R.aluCalc~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Selector11~5_combout\,
	datae => \ALT_INV_R.aluRes\(21),
	dataf => \ALT_INV_R.aluCalc~q\,
	combout => \vAluRes~18_combout\);

-- Location: LABCELL_X80_Y4_N33
\vAluRes~20\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~20_combout\ = ( \Selector9~5_combout\ & ( (\R.aluRes\(23)) # (\R.aluCalc~q\) ) ) # ( !\Selector9~5_combout\ & ( (!\R.aluCalc~q\ & \R.aluRes\(23)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011001100000000001100110000110011111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluCalc~q\,
	datad => \ALT_INV_R.aluRes\(23),
	dataf => \ALT_INV_Selector9~5_combout\,
	combout => \vAluRes~20_combout\);

-- Location: LABCELL_X80_Y4_N24
\vAluRes~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~21_combout\ = (!\R.aluCalc~q\ & (\R.aluRes\(24))) # (\R.aluCalc~q\ & ((\Selector8~4_combout\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000110000111111000011000011111100001100001111110000110000111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluCalc~q\,
	datac => \ALT_INV_R.aluRes\(24),
	datad => \ALT_INV_Selector8~4_combout\,
	combout => \vAluRes~21_combout\);

-- Location: LABCELL_X83_Y3_N36
\vAluRes~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~22_combout\ = ( \R.aluRes\(25) & ( \R.aluCalc~q\ & ( \Selector7~3_combout\ ) ) ) # ( !\R.aluRes\(25) & ( \R.aluCalc~q\ & ( \Selector7~3_combout\ ) ) ) # ( \R.aluRes\(25) & ( !\R.aluCalc~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Selector7~3_combout\,
	datae => \ALT_INV_R.aluRes\(25),
	dataf => \ALT_INV_R.aluCalc~q\,
	combout => \vAluRes~22_combout\);

-- Location: MLABCELL_X78_Y7_N27
\vAluRes~23\ : cyclonev_lcell_comb
-- Equation(s):
-- \vAluRes~23_combout\ = (!\R.aluCalc~q\ & (\R.aluRes\(26))) # (\R.aluCalc~q\ & ((\Selector6~2_combout\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100001111001100110000111100110011000011110011001100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.aluRes\(26),
	datac => \ALT_INV_Selector6~2_combout\,
	datad => \ALT_INV_R.aluCalc~q\,
	combout => \vAluRes~23_combout\);

-- Location: LABCELL_X51_Y2_N24
\Mux221~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux221~1_combout\ = ( \Mux162~0_combout\ & ( \Mux221~0_combout\ ) ) # ( !\Mux162~0_combout\ & ( \Mux221~0_combout\ ) ) # ( \Mux162~0_combout\ & ( !\Mux221~0_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111111111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datae => \ALT_INV_Mux162~0_combout\,
	dataf => \ALT_INV_Mux221~0_combout\,
	combout => \Mux221~1_combout\);

-- Location: LABCELL_X80_Y1_N24
\NxR~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR~6_combout\ = ( \R.ctrlState.Calc~q\ & ( (!\R.curInst\(4) & (\Mux53~1_combout\ & (!\R.curInst\(6) & \R.curInst\(5)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000001000000000000000100000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(4),
	datab => \ALT_INV_Mux53~1_combout\,
	datac => \ALT_INV_R.curInst\(6),
	datad => \ALT_INV_R.curInst\(5),
	dataf => \ALT_INV_R.ctrlState.Calc~q\,
	combout => \NxR~6_combout\);

-- Location: FF_X80_Y1_N25
\R.memWrite\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR~6_combout\,
	asdata => \~GND~combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sclr => \R.ctrlState.Fetch~q\,
	sload => \R.ctrlState.ReadReg~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.memWrite~q\);

-- Location: LABCELL_X66_Y1_N48
\Mux194~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux194~0_combout\ = ( \R.curInst\(14) & ( \Mux114~13_combout\ & ( (!\R.curInst\(13) & ((\Mux122~13_combout\) # (\R.curInst\(12)))) ) ) ) # ( !\R.curInst\(14) & ( \Mux114~13_combout\ & ( (!\R.curInst\(12) & ((!\R.curInst\(13) & (\Mux122~13_combout\)) # 
-- (\R.curInst\(13) & ((\Mux98~13_combout\))))) # (\R.curInst\(12) & (((!\R.curInst\(13))))) ) ) ) # ( \R.curInst\(14) & ( !\Mux114~13_combout\ & ( (!\R.curInst\(12) & (\Mux122~13_combout\ & !\R.curInst\(13))) ) ) ) # ( !\R.curInst\(14) & ( 
-- !\Mux114~13_combout\ & ( (!\R.curInst\(12) & ((!\R.curInst\(13) & (\Mux122~13_combout\)) # (\R.curInst\(13) & ((\Mux98~13_combout\))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010001000001010001000100000000001110111000010100111011100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(12),
	datab => \ALT_INV_Mux122~13_combout\,
	datac => \ALT_INV_Mux98~13_combout\,
	datad => \ALT_INV_R.curInst\(13),
	datae => \ALT_INV_R.curInst\(14),
	dataf => \ALT_INV_Mux114~13_combout\,
	combout => \Mux194~0_combout\);

-- Location: MLABCELL_X59_Y4_N0
\Mux193~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux193~0_combout\ = ( \R.curInst\(12) & ( \Mux113~13_combout\ & ( !\R.curInst\(13) ) ) ) # ( !\R.curInst\(12) & ( \Mux113~13_combout\ & ( (!\R.curInst\(13) & (((\Mux121~13_combout\)))) # (\R.curInst\(13) & (\Mux97~13_combout\ & ((!\R.curInst\(14))))) ) ) 
-- ) # ( !\R.curInst\(12) & ( !\Mux113~13_combout\ & ( (!\R.curInst\(13) & (((\Mux121~13_combout\)))) # (\R.curInst\(13) & (\Mux97~13_combout\ & ((!\R.curInst\(14))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011010100110000000000000000000000110101001100001111000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux97~13_combout\,
	datab => \ALT_INV_Mux121~13_combout\,
	datac => \ALT_INV_R.curInst\(13),
	datad => \ALT_INV_R.curInst\(14),
	datae => \ALT_INV_R.curInst\(12),
	dataf => \ALT_INV_Mux113~13_combout\,
	combout => \Mux193~0_combout\);

-- Location: MLABCELL_X59_Y4_N45
\Mux192~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux192~0_combout\ = ( \R.curInst\(12) & ( \Mux120~13_combout\ & ( (\Mux112~13_combout\ & !\R.curInst\(13)) ) ) ) # ( !\R.curInst\(12) & ( \Mux120~13_combout\ & ( (!\R.curInst\(13)) # ((\Mux96~13_combout\ & !\R.curInst\(14))) ) ) ) # ( \R.curInst\(12) & ( 
-- !\Mux120~13_combout\ & ( (\Mux112~13_combout\ & !\R.curInst\(13)) ) ) ) # ( !\R.curInst\(12) & ( !\Mux120~13_combout\ & ( (\Mux96~13_combout\ & (!\R.curInst\(14) & \R.curInst\(13))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001000100000011110000000011111111010001000000111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux96~13_combout\,
	datab => \ALT_INV_R.curInst\(14),
	datac => \ALT_INV_Mux112~13_combout\,
	datad => \ALT_INV_R.curInst\(13),
	datae => \ALT_INV_R.curInst\(12),
	dataf => \ALT_INV_Mux120~13_combout\,
	combout => \Mux192~0_combout\);

-- Location: LABCELL_X60_Y4_N48
\Mux191~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux191~0_combout\ = ( \Mux111~13_combout\ & ( \R.curInst\(12) & ( !\R.curInst\(13) ) ) ) # ( \Mux111~13_combout\ & ( !\R.curInst\(12) & ( (!\R.curInst\(13) & (\Mux119~13_combout\)) # (\R.curInst\(13) & (((!\R.curInst\(14) & \Mux95~13_combout\)))) ) ) ) # 
-- ( !\Mux111~13_combout\ & ( !\R.curInst\(12) & ( (!\R.curInst\(13) & (\Mux119~13_combout\)) # (\R.curInst\(13) & (((!\R.curInst\(14) & \Mux95~13_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010100001100010101010000110000000000000000001111111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux119~13_combout\,
	datab => \ALT_INV_R.curInst\(14),
	datac => \ALT_INV_Mux95~13_combout\,
	datad => \ALT_INV_R.curInst\(13),
	datae => \ALT_INV_Mux111~13_combout\,
	dataf => \ALT_INV_R.curInst\(12),
	combout => \Mux191~0_combout\);

-- Location: LABCELL_X74_Y4_N24
\Mux190~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux190~0_combout\ = ( \Mux94~13_combout\ & ( \Mux118~13_combout\ & ( (!\R.curInst\(12) & ((!\R.curInst\(13)) # ((!\R.curInst\(14))))) # (\R.curInst\(12) & (!\R.curInst\(13) & ((\Mux110~13_combout\)))) ) ) ) # ( !\Mux94~13_combout\ & ( \Mux118~13_combout\ 
-- & ( (!\R.curInst\(13) & ((!\R.curInst\(12)) # (\Mux110~13_combout\))) ) ) ) # ( \Mux94~13_combout\ & ( !\Mux118~13_combout\ & ( (!\R.curInst\(12) & (\R.curInst\(13) & (!\R.curInst\(14)))) # (\R.curInst\(12) & (!\R.curInst\(13) & ((\Mux110~13_combout\)))) 
-- ) ) ) # ( !\Mux94~13_combout\ & ( !\Mux118~13_combout\ & ( (\R.curInst\(12) & (!\R.curInst\(13) & \Mux110~13_combout\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001000100001000000110010010001000110011001010100011101100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(12),
	datab => \ALT_INV_R.curInst\(13),
	datac => \ALT_INV_R.curInst\(14),
	datad => \ALT_INV_Mux110~13_combout\,
	datae => \ALT_INV_Mux94~13_combout\,
	dataf => \ALT_INV_Mux118~13_combout\,
	combout => \Mux190~0_combout\);

-- Location: MLABCELL_X59_Y4_N36
\Mux189~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux189~0_combout\ = ( \R.curInst\(13) & ( \Mux93~13_combout\ & ( (!\R.curInst\(12) & !\R.curInst\(14)) ) ) ) # ( !\R.curInst\(13) & ( \Mux93~13_combout\ & ( (!\R.curInst\(12) & ((\Mux117~13_combout\))) # (\R.curInst\(12) & (\Mux109~13_combout\)) ) ) ) # 
-- ( !\R.curInst\(13) & ( !\Mux93~13_combout\ & ( (!\R.curInst\(12) & ((\Mux117~13_combout\))) # (\R.curInst\(12) & (\Mux109~13_combout\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001101100011011000000000000000000011011000110111010101000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(12),
	datab => \ALT_INV_Mux109~13_combout\,
	datac => \ALT_INV_Mux117~13_combout\,
	datad => \ALT_INV_R.curInst\(14),
	datae => \ALT_INV_R.curInst\(13),
	dataf => \ALT_INV_Mux93~13_combout\,
	combout => \Mux189~0_combout\);

-- Location: MLABCELL_X59_Y4_N6
\Mux188~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux188~0_combout\ = ( \R.curInst\(12) & ( \Mux116~13_combout\ & ( (!\R.curInst\(13) & \Mux108~13_combout\) ) ) ) # ( !\R.curInst\(12) & ( \Mux116~13_combout\ & ( (!\R.curInst\(13)) # ((!\R.curInst\(14) & \Mux92~13_combout\)) ) ) ) # ( \R.curInst\(12) & ( 
-- !\Mux116~13_combout\ & ( (!\R.curInst\(13) & \Mux108~13_combout\) ) ) ) # ( !\R.curInst\(12) & ( !\Mux116~13_combout\ & ( (\R.curInst\(13) & (!\R.curInst\(14) & \Mux92~13_combout\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010000000100000000001010101010101110101011100000000010101010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(13),
	datab => \ALT_INV_R.curInst\(14),
	datac => \ALT_INV_Mux92~13_combout\,
	datad => \ALT_INV_Mux108~13_combout\,
	datae => \ALT_INV_R.curInst\(12),
	dataf => \ALT_INV_Mux116~13_combout\,
	combout => \Mux188~0_combout\);

-- Location: MLABCELL_X59_Y4_N18
\Mux187~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux187~0_combout\ = ( \R.curInst\(12) & ( \Mux115~13_combout\ & ( (!\R.curInst\(13) & \Mux107~13_combout\) ) ) ) # ( !\R.curInst\(12) & ( \Mux115~13_combout\ & ( (!\R.curInst\(13)) # ((\Mux91~13_combout\ & !\R.curInst\(14))) ) ) ) # ( \R.curInst\(12) & ( 
-- !\Mux115~13_combout\ & ( (!\R.curInst\(13) & \Mux107~13_combout\) ) ) ) # ( !\R.curInst\(12) & ( !\Mux115~13_combout\ & ( (\R.curInst\(13) & (\Mux91~13_combout\ & !\R.curInst\(14))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000000001000100010001010101111101010100010001000100010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(13),
	datab => \ALT_INV_Mux107~13_combout\,
	datac => \ALT_INV_Mux91~13_combout\,
	datad => \ALT_INV_R.curInst\(14),
	datae => \ALT_INV_R.curInst\(12),
	dataf => \ALT_INV_Mux115~13_combout\,
	combout => \Mux187~0_combout\);

-- Location: LABCELL_X71_Y1_N51
\Mux202~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux202~0_combout\ = ( \Mux122~13_combout\ & ( (!\R.curInst\(13) & (((\R.curInst\(12))))) # (\R.curInst\(13) & (!\R.curInst\(14) & (!\R.curInst\(12) & \Mux106~13_combout\))) ) ) # ( !\Mux122~13_combout\ & ( (!\R.curInst\(14) & (\R.curInst\(13) & 
-- (!\R.curInst\(12) & \Mux106~13_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000100000000011000010110000000000001000000000110000101100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(14),
	datab => \ALT_INV_R.curInst\(13),
	datac => \ALT_INV_R.curInst\(12),
	datad => \ALT_INV_Mux106~13_combout\,
	datae => \ALT_INV_Mux122~13_combout\,
	combout => \Mux202~0_combout\);

-- Location: MLABCELL_X59_Y4_N51
\Mux201~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux201~0_combout\ = ( \Mux105~13_combout\ & ( (!\R.curInst\(12) & (!\R.curInst\(14) & ((\R.curInst\(13))))) # (\R.curInst\(12) & (((\Mux121~13_combout\ & !\R.curInst\(13))))) ) ) # ( !\Mux105~13_combout\ & ( (\R.curInst\(12) & (\Mux121~13_combout\ & 
-- !\R.curInst\(13))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000000000001010000000000000101100010000000010110001000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(12),
	datab => \ALT_INV_R.curInst\(14),
	datac => \ALT_INV_Mux121~13_combout\,
	datad => \ALT_INV_R.curInst\(13),
	dataf => \ALT_INV_Mux105~13_combout\,
	combout => \Mux201~0_combout\);

-- Location: MLABCELL_X59_Y4_N54
\Mux200~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux200~0_combout\ = ( \R.curInst\(13) & ( \Mux120~13_combout\ & ( (!\R.curInst\(12) & (\Mux104~13_combout\ & !\R.curInst\(14))) ) ) ) # ( !\R.curInst\(13) & ( \Mux120~13_combout\ & ( \R.curInst\(12) ) ) ) # ( \R.curInst\(13) & ( !\Mux120~13_combout\ & ( 
-- (!\R.curInst\(12) & (\Mux104~13_combout\ & !\R.curInst\(14))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011000000000000110011001100110000110000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_R.curInst\(12),
	datac => \ALT_INV_Mux104~13_combout\,
	datad => \ALT_INV_R.curInst\(14),
	datae => \ALT_INV_R.curInst\(13),
	dataf => \ALT_INV_Mux120~13_combout\,
	combout => \Mux200~0_combout\);

-- Location: LABCELL_X71_Y1_N9
\Mux199~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux199~0_combout\ = ( \Mux103~13_combout\ & ( \R.curInst\(12) & ( (!\R.curInst\(13) & \Mux119~13_combout\) ) ) ) # ( !\Mux103~13_combout\ & ( \R.curInst\(12) & ( (!\R.curInst\(13) & \Mux119~13_combout\) ) ) ) # ( \Mux103~13_combout\ & ( !\R.curInst\(12) 
-- & ( (!\R.curInst\(14) & \R.curInst\(13)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000001000100010001000001100000011000000110000001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(14),
	datab => \ALT_INV_R.curInst\(13),
	datac => \ALT_INV_Mux119~13_combout\,
	datae => \ALT_INV_Mux103~13_combout\,
	dataf => \ALT_INV_R.curInst\(12),
	combout => \Mux199~0_combout\);

-- Location: MLABCELL_X59_Y4_N48
\Mux198~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux198~0_combout\ = ( \Mux118~13_combout\ & ( (!\R.curInst\(12) & (!\R.curInst\(14) & (\Mux102~13_combout\ & \R.curInst\(13)))) # (\R.curInst\(12) & (((!\R.curInst\(13))))) ) ) # ( !\Mux118~13_combout\ & ( (!\R.curInst\(12) & (!\R.curInst\(14) & 
-- (\Mux102~13_combout\ & \R.curInst\(13)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000001000000000000000100001010101000010000101010100001000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(12),
	datab => \ALT_INV_R.curInst\(14),
	datac => \ALT_INV_Mux102~13_combout\,
	datad => \ALT_INV_R.curInst\(13),
	dataf => \ALT_INV_Mux118~13_combout\,
	combout => \Mux198~0_combout\);

-- Location: MLABCELL_X59_Y4_N24
\Mux197~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux197~0_combout\ = ( \R.curInst\(13) & ( \Mux117~13_combout\ & ( (\Mux101~13_combout\ & (!\R.curInst\(14) & !\R.curInst\(12))) ) ) ) # ( !\R.curInst\(13) & ( \Mux117~13_combout\ & ( \R.curInst\(12) ) ) ) # ( \R.curInst\(13) & ( !\Mux117~13_combout\ & ( 
-- (\Mux101~13_combout\ & (!\R.curInst\(14) & !\R.curInst\(12))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010001000000000000000000111111110100010000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux101~13_combout\,
	datab => \ALT_INV_R.curInst\(14),
	datad => \ALT_INV_R.curInst\(12),
	datae => \ALT_INV_R.curInst\(13),
	dataf => \ALT_INV_Mux117~13_combout\,
	combout => \Mux197~0_combout\);

-- Location: MLABCELL_X59_Y4_N33
\Mux196~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux196~0_combout\ = ( \Mux116~13_combout\ & ( (!\R.curInst\(13) & (((\R.curInst\(12))))) # (\R.curInst\(13) & (!\R.curInst\(14) & (\Mux100~13_combout\ & !\R.curInst\(12)))) ) ) # ( !\Mux116~13_combout\ & ( (\R.curInst\(13) & (!\R.curInst\(14) & 
-- (\Mux100~13_combout\ & !\R.curInst\(12)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010000000000000001000000000000000100101010100000010010101010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(13),
	datab => \ALT_INV_R.curInst\(14),
	datac => \ALT_INV_Mux100~13_combout\,
	datad => \ALT_INV_R.curInst\(12),
	dataf => \ALT_INV_Mux116~13_combout\,
	combout => \Mux196~0_combout\);

-- Location: MLABCELL_X59_Y4_N30
\Mux195~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux195~0_combout\ = ( \Mux115~13_combout\ & ( (!\R.curInst\(13) & (((\R.curInst\(12))))) # (\R.curInst\(13) & (!\R.curInst\(14) & (!\R.curInst\(12) & \Mux99~13_combout\))) ) ) # ( !\Mux115~13_combout\ & ( (\R.curInst\(13) & (!\R.curInst\(14) & 
-- (!\R.curInst\(12) & \Mux99~13_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001000000000000000100000000001010010010100000101001001010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(13),
	datab => \ALT_INV_R.curInst\(14),
	datac => \ALT_INV_R.curInst\(12),
	datad => \ALT_INV_Mux99~13_combout\,
	dataf => \ALT_INV_Mux115~13_combout\,
	combout => \Mux195~0_combout\);

-- Location: LABCELL_X30_Y1_N39
\Mux210~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux210~0_combout\ = ( \Mux221~0_combout\ & ( \Mux114~13_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Mux114~13_combout\,
	dataf => \ALT_INV_Mux221~0_combout\,
	combout => \Mux210~0_combout\);

-- Location: LABCELL_X51_Y4_N48
\Mux209~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux209~0_combout\ = ( \Mux221~0_combout\ & ( \Mux113~13_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000110011001100110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Mux113~13_combout\,
	dataf => \ALT_INV_Mux221~0_combout\,
	combout => \Mux209~0_combout\);

-- Location: LABCELL_X51_Y4_N57
\Mux208~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux208~0_combout\ = ( \Mux112~13_combout\ & ( \Mux221~0_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000001010101010101010101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux221~0_combout\,
	dataf => \ALT_INV_Mux112~13_combout\,
	combout => \Mux208~0_combout\);

-- Location: LABCELL_X30_Y1_N30
\Mux207~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux207~0_combout\ = ( \Mux221~0_combout\ & ( \Mux111~13_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000110011001100110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Mux111~13_combout\,
	dataf => \ALT_INV_Mux221~0_combout\,
	combout => \Mux207~0_combout\);

-- Location: LABCELL_X51_Y4_N24
\Mux206~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux206~0_combout\ = ( \Mux110~13_combout\ & ( \Mux221~0_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Mux221~0_combout\,
	dataf => \ALT_INV_Mux110~13_combout\,
	combout => \Mux206~0_combout\);

-- Location: LABCELL_X51_Y2_N30
\Mux205~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux205~0_combout\ = ( \Mux221~0_combout\ & ( \Mux109~13_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Mux109~13_combout\,
	dataf => \ALT_INV_Mux221~0_combout\,
	combout => \Mux205~0_combout\);

-- Location: LABCELL_X51_Y4_N6
\Mux204~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux204~0_combout\ = ( \Mux108~13_combout\ & ( \Mux221~0_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Mux221~0_combout\,
	dataf => \ALT_INV_Mux108~13_combout\,
	combout => \Mux204~0_combout\);

-- Location: MLABCELL_X59_Y4_N15
\Mux203~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux203~0_combout\ = ( \Mux221~0_combout\ & ( \Mux107~13_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Mux107~13_combout\,
	datae => \ALT_INV_Mux221~0_combout\,
	combout => \Mux203~0_combout\);

-- Location: LABCELL_X51_Y2_N48
\Mux218~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux218~0_combout\ = ( \Mux221~0_combout\ & ( \Mux122~13_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Mux122~13_combout\,
	dataf => \ALT_INV_Mux221~0_combout\,
	combout => \Mux218~0_combout\);

-- Location: LABCELL_X83_Y4_N45
\Mux217~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux217~0_combout\ = ( \Mux121~13_combout\ & ( \Mux221~0_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Mux221~0_combout\,
	dataf => \ALT_INV_Mux121~13_combout\,
	combout => \Mux217~0_combout\);

-- Location: LABCELL_X71_Y5_N54
\Mux216~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux216~0_combout\ = ( \Mux221~0_combout\ & ( \Mux120~13_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000110011001100110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Mux120~13_combout\,
	dataf => \ALT_INV_Mux221~0_combout\,
	combout => \Mux216~0_combout\);

-- Location: LABCELL_X51_Y4_N12
\Mux215~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux215~0_combout\ = ( \Mux119~13_combout\ & ( \Mux221~0_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Mux221~0_combout\,
	dataf => \ALT_INV_Mux119~13_combout\,
	combout => \Mux215~0_combout\);

-- Location: LABCELL_X51_Y4_N42
\Mux214~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux214~0_combout\ = ( \Mux118~13_combout\ & ( \Mux221~0_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ALT_INV_Mux221~0_combout\,
	dataf => \ALT_INV_Mux118~13_combout\,
	combout => \Mux214~0_combout\);

-- Location: MLABCELL_X52_Y5_N39
\Mux213~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux213~0_combout\ = ( \Mux221~0_combout\ & ( \Mux117~13_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000001010101010101010101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux117~13_combout\,
	dataf => \ALT_INV_Mux221~0_combout\,
	combout => \Mux213~0_combout\);

-- Location: LABCELL_X51_Y4_N36
\Mux212~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux212~0_combout\ = ( \Mux221~0_combout\ & ( \Mux116~13_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000110011001100110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ALT_INV_Mux116~13_combout\,
	dataf => \ALT_INV_Mux221~0_combout\,
	combout => \Mux212~0_combout\);

-- Location: MLABCELL_X52_Y5_N33
\Mux211~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Mux211~0_combout\ = ( \Mux221~0_combout\ & ( \Mux115~13_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000001010101010101010101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_Mux115~13_combout\,
	dataf => \ALT_INV_Mux221~0_combout\,
	combout => \Mux211~0_combout\);

-- Location: LABCELL_X80_Y1_N42
\NxR~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \NxR~7_combout\ = ( \Mux53~1_combout\ & ( (!\R.curInst\(4) & (\R.ctrlState.Calc~q\ & \Mux154~0_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000010000000100000001000000010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_R.curInst\(4),
	datab => \ALT_INV_R.ctrlState.Calc~q\,
	datac => \ALT_INV_Mux154~0_combout\,
	dataf => \ALT_INV_Mux53~1_combout\,
	combout => \NxR~7_combout\);

-- Location: FF_X80_Y1_N43
\R.memRead\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \csi_clk~inputCLKENA0_outclk\,
	d => \NxR~7_combout\,
	asdata => \~GND~combout\,
	clrn => \rsi_reset_n~inputCLKENA0_outclk\,
	sclr => \R.ctrlState.Fetch~q\,
	sload => \R.ctrlState.ReadReg~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \R.memRead~q\);

-- Location: IOIBUF_X8_Y81_N35
\avm_i_waitrequest~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_i_waitrequest,
	o => \avm_i_waitrequest~input_o\);

-- Location: IOIBUF_X30_Y81_N52
\avm_d_waitrequest~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_avm_d_waitrequest,
	o => \avm_d_waitrequest~input_o\);
END structure;


