-- riscv_simulation.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity riscv_simulation is
	port (
		leds_export : out std_logic_vector(7 downto 0)   -- leds.export
	);
end entity riscv_simulation;

architecture rtl of riscv_simulation is
	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component riscv_simulation_onchip_memory2_0 is
		port (
			address     : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			address2    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk         : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			freeze      : in  std_logic                     := 'X'              -- freeze
		);
	end component riscv_simulation_onchip_memory2_0;

	component riscv_simulation_pio_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component riscv_simulation_pio_0;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	component Core is
		port (
			csi_clk           : in  std_logic                     := 'X';             -- clk
			avm_d_address     : out std_logic_vector(31 downto 0);                    -- address
			avm_d_byteenable  : out std_logic_vector(3 downto 0);                     -- byteenable
			avm_d_write       : out std_logic;                                        -- write
			avm_d_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			avm_d_read        : out std_logic;                                        -- read
			avm_d_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			avm_d_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			avm_i_address     : out std_logic_vector(31 downto 0);                    -- address
			avm_i_read        : out std_logic;                                        -- read
			avm_i_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			avm_i_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			rsi_reset_n       : in  std_logic                     := 'X'              -- reset_n
		);
	end component Core;

	component riscv_simulation_mm_interconnect_0 is
		port (
			clock_source_0_clk_clk                            : in  std_logic                     := 'X';             -- clk
			rv32ui_fsmd_0_reset_n_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			rv32ui_fsmd_0_data_address                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			rv32ui_fsmd_0_data_waitrequest                    : out std_logic;                                        -- waitrequest
			rv32ui_fsmd_0_data_byteenable                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			rv32ui_fsmd_0_data_read                           : in  std_logic                     := 'X';             -- read
			rv32ui_fsmd_0_data_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			rv32ui_fsmd_0_data_write                          : in  std_logic                     := 'X';             -- write
			rv32ui_fsmd_0_data_writedata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			onchip_memory2_0_s2_address                       : out std_logic_vector(12 downto 0);                    -- address
			onchip_memory2_0_s2_write                         : out std_logic;                                        -- write
			onchip_memory2_0_s2_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s2_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s2_byteenable                    : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s2_chipselect                    : out std_logic;                                        -- chipselect
			onchip_memory2_0_s2_clken                         : out std_logic;                                        -- clken
			pio_0_s1_address                                  : out std_logic_vector(1 downto 0);                     -- address
			pio_0_s1_write                                    : out std_logic;                                        -- write
			pio_0_s1_readdata                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_0_s1_writedata                                : out std_logic_vector(31 downto 0);                    -- writedata
			pio_0_s1_chipselect                               : out std_logic                                         -- chipselect
		);
	end component riscv_simulation_mm_interconnect_0;

	component riscv_simulation_mm_interconnect_1 is
		port (
			clock_source_0_clk_clk                            : in  std_logic                     := 'X';             -- clk
			rv32ui_fsmd_0_reset_n_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			rv32ui_fsmd_0_instruction_address                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			rv32ui_fsmd_0_instruction_waitrequest             : out std_logic;                                        -- waitrequest
			rv32ui_fsmd_0_instruction_read                    : in  std_logic                     := 'X';             -- read
			rv32ui_fsmd_0_instruction_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			onchip_memory2_0_s1_address                       : out std_logic_vector(12 downto 0);                    -- address
			onchip_memory2_0_s1_write                         : out std_logic;                                        -- write
			onchip_memory2_0_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                    : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                    : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_clken                         : out std_logic                                         -- clken
		);
	end component riscv_simulation_mm_interconnect_1;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal clock_source_0_clk_clk                           : std_logic;                     -- clock_source_0:clk -> [mm_interconnect_0:clock_source_0_clk_clk, mm_interconnect_1:clock_source_0_clk_clk, onchip_memory2_0:clk, pio_0:clk, reset_source_0:clk, rst_controller:clk, rv32ui_fsmd_0:csi_clk]
	signal rv32ui_fsmd_0_data_readdata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:rv32ui_fsmd_0_data_readdata -> rv32ui_fsmd_0:avm_d_readdata
	signal rv32ui_fsmd_0_data_waitrequest                   : std_logic;                     -- mm_interconnect_0:rv32ui_fsmd_0_data_waitrequest -> rv32ui_fsmd_0:avm_d_waitrequest
	signal rv32ui_fsmd_0_data_address                       : std_logic_vector(31 downto 0); -- rv32ui_fsmd_0:avm_d_address -> mm_interconnect_0:rv32ui_fsmd_0_data_address
	signal rv32ui_fsmd_0_data_byteenable                    : std_logic_vector(3 downto 0);  -- rv32ui_fsmd_0:avm_d_byteenable -> mm_interconnect_0:rv32ui_fsmd_0_data_byteenable
	signal rv32ui_fsmd_0_data_read                          : std_logic;                     -- rv32ui_fsmd_0:avm_d_read -> mm_interconnect_0:rv32ui_fsmd_0_data_read
	signal rv32ui_fsmd_0_data_write                         : std_logic;                     -- rv32ui_fsmd_0:avm_d_write -> mm_interconnect_0:rv32ui_fsmd_0_data_write
	signal rv32ui_fsmd_0_data_writedata                     : std_logic_vector(31 downto 0); -- rv32ui_fsmd_0:avm_d_writedata -> mm_interconnect_0:rv32ui_fsmd_0_data_writedata
	signal mm_interconnect_0_pio_0_s1_chipselect            : std_logic;                     -- mm_interconnect_0:pio_0_s1_chipselect -> pio_0:chipselect
	signal mm_interconnect_0_pio_0_s1_readdata              : std_logic_vector(31 downto 0); -- pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	signal mm_interconnect_0_pio_0_s1_address               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_0_s1_address -> pio_0:address
	signal mm_interconnect_0_pio_0_s1_write                 : std_logic;                     -- mm_interconnect_0:pio_0_s1_write -> mm_interconnect_0_pio_0_s1_write:in
	signal mm_interconnect_0_pio_0_s1_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_0_s1_writedata -> pio_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s2_chipselect : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s2_chipselect -> onchip_memory2_0:chipselect2
	signal mm_interconnect_0_onchip_memory2_0_s2_readdata   : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata2 -> mm_interconnect_0:onchip_memory2_0_s2_readdata
	signal mm_interconnect_0_onchip_memory2_0_s2_address    : std_logic_vector(12 downto 0); -- mm_interconnect_0:onchip_memory2_0_s2_address -> onchip_memory2_0:address2
	signal mm_interconnect_0_onchip_memory2_0_s2_byteenable : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s2_byteenable -> onchip_memory2_0:byteenable2
	signal mm_interconnect_0_onchip_memory2_0_s2_write      : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s2_write -> onchip_memory2_0:write2
	signal mm_interconnect_0_onchip_memory2_0_s2_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_0_s2_writedata -> onchip_memory2_0:writedata2
	signal mm_interconnect_0_onchip_memory2_0_s2_clken      : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s2_clken -> onchip_memory2_0:clken2
	signal rv32ui_fsmd_0_instruction_readdata               : std_logic_vector(31 downto 0); -- mm_interconnect_1:rv32ui_fsmd_0_instruction_readdata -> rv32ui_fsmd_0:avm_i_readdata
	signal rv32ui_fsmd_0_instruction_waitrequest            : std_logic;                     -- mm_interconnect_1:rv32ui_fsmd_0_instruction_waitrequest -> rv32ui_fsmd_0:avm_i_waitrequest
	signal rv32ui_fsmd_0_instruction_address                : std_logic_vector(31 downto 0); -- rv32ui_fsmd_0:avm_i_address -> mm_interconnect_1:rv32ui_fsmd_0_instruction_address
	signal rv32ui_fsmd_0_instruction_read                   : std_logic;                     -- rv32ui_fsmd_0:avm_i_read -> mm_interconnect_1:rv32ui_fsmd_0_instruction_read
	signal mm_interconnect_1_onchip_memory2_0_s1_chipselect : std_logic;                     -- mm_interconnect_1:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_1_onchip_memory2_0_s1_readdata   : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata -> mm_interconnect_1:onchip_memory2_0_s1_readdata
	signal mm_interconnect_1_onchip_memory2_0_s1_address    : std_logic_vector(12 downto 0); -- mm_interconnect_1:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_1_onchip_memory2_0_s1_byteenable : std_logic_vector(3 downto 0);  -- mm_interconnect_1:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_1_onchip_memory2_0_s1_write      : std_logic;                     -- mm_interconnect_1:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_1_onchip_memory2_0_s1_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_1:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_1_onchip_memory2_0_s1_clken      : std_logic;                     -- mm_interconnect_1:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal rst_controller_reset_out_reset                   : std_logic;                     -- rst_controller:reset_out -> [mm_interconnect_0:rv32ui_fsmd_0_reset_n_reset_bridge_in_reset_reset, mm_interconnect_1:rv32ui_fsmd_0_reset_n_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req               : std_logic;                     -- rst_controller:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	signal reset_source_0_reset_reset                       : std_logic;                     -- reset_source_0:reset -> rst_controller:reset_in0
	signal mm_interconnect_0_pio_0_s1_write_ports_inv       : std_logic;                     -- mm_interconnect_0_pio_0_s1_write:inv -> pio_0:write_n
	signal rst_controller_reset_out_reset_ports_inv         : std_logic;                     -- rst_controller_reset_out_reset:inv -> [pio_0:reset_n, rv32ui_fsmd_0:rsi_reset_n]

begin

	clock_source_0 : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50,
			CLOCK_UNIT => 1000000
		)
		port map (
			clk => clock_source_0_clk_clk  -- clk.clk
		);

	onchip_memory2_0 : component riscv_simulation_onchip_memory2_0
		port map (
			address     => mm_interconnect_1_onchip_memory2_0_s1_address,    --     s1.address
			clken       => mm_interconnect_1_onchip_memory2_0_s1_clken,      --       .clken
			chipselect  => mm_interconnect_1_onchip_memory2_0_s1_chipselect, --       .chipselect
			write       => mm_interconnect_1_onchip_memory2_0_s1_write,      --       .write
			readdata    => mm_interconnect_1_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_1_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_1_onchip_memory2_0_s1_byteenable, --       .byteenable
			address2    => mm_interconnect_0_onchip_memory2_0_s2_address,    --     s2.address
			chipselect2 => mm_interconnect_0_onchip_memory2_0_s2_chipselect, --       .chipselect
			clken2      => mm_interconnect_0_onchip_memory2_0_s2_clken,      --       .clken
			write2      => mm_interconnect_0_onchip_memory2_0_s2_write,      --       .write
			readdata2   => mm_interconnect_0_onchip_memory2_0_s2_readdata,   --       .readdata
			writedata2  => mm_interconnect_0_onchip_memory2_0_s2_writedata,  --       .writedata
			byteenable2 => mm_interconnect_0_onchip_memory2_0_s2_byteenable, --       .byteenable
			clk         => clock_source_0_clk_clk,                           --   clk1.clk
			reset       => rst_controller_reset_out_reset,                   -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,               --       .reset_req
			freeze      => '0'                                               -- (terminated)
		);

	pio_0 : component riscv_simulation_pio_0
		port map (
			clk        => clock_source_0_clk_clk,                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_pio_0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_0_s1_readdata,        --                    .readdata
			out_port   => leds_export                                 -- external_connection.export
		);

	reset_source_0 : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 1,
			INITIAL_RESET_CYCLES => 10
		)
		port map (
			reset => reset_source_0_reset_reset, -- reset.reset
			clk   => clock_source_0_clk_clk      --   clk.clk
		);

	rv32ui_fsmd_0 : component Core
		port map (
			csi_clk           => clock_source_0_clk_clk,                   --       clock.clk
			avm_d_address     => rv32ui_fsmd_0_data_address,               --        data.address
			avm_d_byteenable  => rv32ui_fsmd_0_data_byteenable,            --            .byteenable
			avm_d_write       => rv32ui_fsmd_0_data_write,                 --            .write
			avm_d_writedata   => rv32ui_fsmd_0_data_writedata,             --            .writedata
			avm_d_read        => rv32ui_fsmd_0_data_read,                  --            .read
			avm_d_readdata    => rv32ui_fsmd_0_data_readdata,              --            .readdata
			avm_d_waitrequest => rv32ui_fsmd_0_data_waitrequest,           --            .waitrequest
			avm_i_address     => rv32ui_fsmd_0_instruction_address,        -- instruction.address
			avm_i_read        => rv32ui_fsmd_0_instruction_read,           --            .read
			avm_i_readdata    => rv32ui_fsmd_0_instruction_readdata,       --            .readdata
			avm_i_waitrequest => rv32ui_fsmd_0_instruction_waitrequest,    --            .waitrequest
			rsi_reset_n       => rst_controller_reset_out_reset_ports_inv  --     reset_n.reset_n
		);

	mm_interconnect_0 : component riscv_simulation_mm_interconnect_0
		port map (
			clock_source_0_clk_clk                            => clock_source_0_clk_clk,                           --                          clock_source_0_clk.clk
			rv32ui_fsmd_0_reset_n_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                   -- rv32ui_fsmd_0_reset_n_reset_bridge_in_reset.reset
			rv32ui_fsmd_0_data_address                        => rv32ui_fsmd_0_data_address,                       --                          rv32ui_fsmd_0_data.address
			rv32ui_fsmd_0_data_waitrequest                    => rv32ui_fsmd_0_data_waitrequest,                   --                                            .waitrequest
			rv32ui_fsmd_0_data_byteenable                     => rv32ui_fsmd_0_data_byteenable,                    --                                            .byteenable
			rv32ui_fsmd_0_data_read                           => rv32ui_fsmd_0_data_read,                          --                                            .read
			rv32ui_fsmd_0_data_readdata                       => rv32ui_fsmd_0_data_readdata,                      --                                            .readdata
			rv32ui_fsmd_0_data_write                          => rv32ui_fsmd_0_data_write,                         --                                            .write
			rv32ui_fsmd_0_data_writedata                      => rv32ui_fsmd_0_data_writedata,                     --                                            .writedata
			onchip_memory2_0_s2_address                       => mm_interconnect_0_onchip_memory2_0_s2_address,    --                         onchip_memory2_0_s2.address
			onchip_memory2_0_s2_write                         => mm_interconnect_0_onchip_memory2_0_s2_write,      --                                            .write
			onchip_memory2_0_s2_readdata                      => mm_interconnect_0_onchip_memory2_0_s2_readdata,   --                                            .readdata
			onchip_memory2_0_s2_writedata                     => mm_interconnect_0_onchip_memory2_0_s2_writedata,  --                                            .writedata
			onchip_memory2_0_s2_byteenable                    => mm_interconnect_0_onchip_memory2_0_s2_byteenable, --                                            .byteenable
			onchip_memory2_0_s2_chipselect                    => mm_interconnect_0_onchip_memory2_0_s2_chipselect, --                                            .chipselect
			onchip_memory2_0_s2_clken                         => mm_interconnect_0_onchip_memory2_0_s2_clken,      --                                            .clken
			pio_0_s1_address                                  => mm_interconnect_0_pio_0_s1_address,               --                                    pio_0_s1.address
			pio_0_s1_write                                    => mm_interconnect_0_pio_0_s1_write,                 --                                            .write
			pio_0_s1_readdata                                 => mm_interconnect_0_pio_0_s1_readdata,              --                                            .readdata
			pio_0_s1_writedata                                => mm_interconnect_0_pio_0_s1_writedata,             --                                            .writedata
			pio_0_s1_chipselect                               => mm_interconnect_0_pio_0_s1_chipselect             --                                            .chipselect
		);

	mm_interconnect_1 : component riscv_simulation_mm_interconnect_1
		port map (
			clock_source_0_clk_clk                            => clock_source_0_clk_clk,                           --                          clock_source_0_clk.clk
			rv32ui_fsmd_0_reset_n_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                   -- rv32ui_fsmd_0_reset_n_reset_bridge_in_reset.reset
			rv32ui_fsmd_0_instruction_address                 => rv32ui_fsmd_0_instruction_address,                --                   rv32ui_fsmd_0_instruction.address
			rv32ui_fsmd_0_instruction_waitrequest             => rv32ui_fsmd_0_instruction_waitrequest,            --                                            .waitrequest
			rv32ui_fsmd_0_instruction_read                    => rv32ui_fsmd_0_instruction_read,                   --                                            .read
			rv32ui_fsmd_0_instruction_readdata                => rv32ui_fsmd_0_instruction_readdata,               --                                            .readdata
			onchip_memory2_0_s1_address                       => mm_interconnect_1_onchip_memory2_0_s1_address,    --                         onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                         => mm_interconnect_1_onchip_memory2_0_s1_write,      --                                            .write
			onchip_memory2_0_s1_readdata                      => mm_interconnect_1_onchip_memory2_0_s1_readdata,   --                                            .readdata
			onchip_memory2_0_s1_writedata                     => mm_interconnect_1_onchip_memory2_0_s1_writedata,  --                                            .writedata
			onchip_memory2_0_s1_byteenable                    => mm_interconnect_1_onchip_memory2_0_s1_byteenable, --                                            .byteenable
			onchip_memory2_0_s1_chipselect                    => mm_interconnect_1_onchip_memory2_0_s1_chipselect, --                                            .chipselect
			onchip_memory2_0_s1_clken                         => mm_interconnect_1_onchip_memory2_0_s1_clken       --                                            .clken
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_source_0_reset_reset,         -- reset_in0.reset
			clk            => clock_source_0_clk_clk,             --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	mm_interconnect_0_pio_0_s1_write_ports_inv <= not mm_interconnect_0_pio_0_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of riscv_simulation
